module DecodeStage_top;

  wire  clock;
  wire  reset;
  wire  io_redirect;
  wire  io_in_0_ready;
  wire  io_in_0_valid;
  wire [31:0] io_in_0_bits_instr;
  wire  io_in_0_bits_exceptionVec_0;
  wire  io_in_0_bits_exceptionVec_1;
  wire  io_in_0_bits_exceptionVec_2;
  wire  io_in_0_bits_exceptionVec_4;
  wire  io_in_0_bits_exceptionVec_5;
  wire  io_in_0_bits_exceptionVec_6;
  wire  io_in_0_bits_exceptionVec_7;
  wire  io_in_0_bits_exceptionVec_8;
  wire  io_in_0_bits_exceptionVec_9;
  wire  io_in_0_bits_exceptionVec_10;
  wire  io_in_0_bits_exceptionVec_11;
  wire  io_in_0_bits_exceptionVec_12;
  wire  io_in_0_bits_exceptionVec_13;
  wire  io_in_0_bits_exceptionVec_14;
  wire  io_in_0_bits_exceptionVec_15;
  wire  io_in_0_bits_exceptionVec_16;
  wire  io_in_0_bits_exceptionVec_17;
  wire  io_in_0_bits_exceptionVec_18;
  wire  io_in_0_bits_exceptionVec_19;
  wire  io_in_0_bits_exceptionVec_20;
  wire  io_in_0_bits_exceptionVec_21;
  wire  io_in_0_bits_exceptionVec_23;
  wire  io_in_0_bits_isFetchMalAddr;
  wire [3:0] io_in_0_bits_trigger;
  wire  io_in_0_bits_preDecodeInfo_isRVC;
  wire [1:0] io_in_0_bits_preDecodeInfo_brType;
  wire  io_in_0_bits_pred_taken;
  wire  io_in_0_bits_crossPageIPFFix;
  wire  io_in_0_bits_ftqPtr_flag;
  wire [5:0] io_in_0_bits_ftqPtr_value;
  wire [3:0] io_in_0_bits_ftqOffset;
  wire  io_in_0_bits_isLastInFtqEntry;
  wire  io_in_1_ready;
  wire  io_in_1_valid;
  wire [31:0] io_in_1_bits_instr;
  wire  io_in_1_bits_exceptionVec_0;
  wire  io_in_1_bits_exceptionVec_1;
  wire  io_in_1_bits_exceptionVec_2;
  wire  io_in_1_bits_exceptionVec_4;
  wire  io_in_1_bits_exceptionVec_5;
  wire  io_in_1_bits_exceptionVec_6;
  wire  io_in_1_bits_exceptionVec_7;
  wire  io_in_1_bits_exceptionVec_8;
  wire  io_in_1_bits_exceptionVec_9;
  wire  io_in_1_bits_exceptionVec_10;
  wire  io_in_1_bits_exceptionVec_11;
  wire  io_in_1_bits_exceptionVec_12;
  wire  io_in_1_bits_exceptionVec_13;
  wire  io_in_1_bits_exceptionVec_14;
  wire  io_in_1_bits_exceptionVec_15;
  wire  io_in_1_bits_exceptionVec_16;
  wire  io_in_1_bits_exceptionVec_17;
  wire  io_in_1_bits_exceptionVec_18;
  wire  io_in_1_bits_exceptionVec_19;
  wire  io_in_1_bits_exceptionVec_20;
  wire  io_in_1_bits_exceptionVec_21;
  wire  io_in_1_bits_exceptionVec_23;
  wire  io_in_1_bits_isFetchMalAddr;
  wire [3:0] io_in_1_bits_trigger;
  wire  io_in_1_bits_preDecodeInfo_isRVC;
  wire [1:0] io_in_1_bits_preDecodeInfo_brType;
  wire  io_in_1_bits_pred_taken;
  wire  io_in_1_bits_crossPageIPFFix;
  wire  io_in_1_bits_ftqPtr_flag;
  wire [5:0] io_in_1_bits_ftqPtr_value;
  wire [3:0] io_in_1_bits_ftqOffset;
  wire  io_in_1_bits_isLastInFtqEntry;
  wire  io_in_2_ready;
  wire  io_in_2_valid;
  wire [31:0] io_in_2_bits_instr;
  wire  io_in_2_bits_exceptionVec_0;
  wire  io_in_2_bits_exceptionVec_1;
  wire  io_in_2_bits_exceptionVec_2;
  wire  io_in_2_bits_exceptionVec_4;
  wire  io_in_2_bits_exceptionVec_5;
  wire  io_in_2_bits_exceptionVec_6;
  wire  io_in_2_bits_exceptionVec_7;
  wire  io_in_2_bits_exceptionVec_8;
  wire  io_in_2_bits_exceptionVec_9;
  wire  io_in_2_bits_exceptionVec_10;
  wire  io_in_2_bits_exceptionVec_11;
  wire  io_in_2_bits_exceptionVec_12;
  wire  io_in_2_bits_exceptionVec_13;
  wire  io_in_2_bits_exceptionVec_14;
  wire  io_in_2_bits_exceptionVec_15;
  wire  io_in_2_bits_exceptionVec_16;
  wire  io_in_2_bits_exceptionVec_17;
  wire  io_in_2_bits_exceptionVec_18;
  wire  io_in_2_bits_exceptionVec_19;
  wire  io_in_2_bits_exceptionVec_20;
  wire  io_in_2_bits_exceptionVec_21;
  wire  io_in_2_bits_exceptionVec_23;
  wire  io_in_2_bits_isFetchMalAddr;
  wire [3:0] io_in_2_bits_trigger;
  wire  io_in_2_bits_preDecodeInfo_isRVC;
  wire [1:0] io_in_2_bits_preDecodeInfo_brType;
  wire  io_in_2_bits_pred_taken;
  wire  io_in_2_bits_crossPageIPFFix;
  wire  io_in_2_bits_ftqPtr_flag;
  wire [5:0] io_in_2_bits_ftqPtr_value;
  wire [3:0] io_in_2_bits_ftqOffset;
  wire  io_in_2_bits_isLastInFtqEntry;
  wire  io_in_3_ready;
  wire  io_in_3_valid;
  wire [31:0] io_in_3_bits_instr;
  wire  io_in_3_bits_exceptionVec_0;
  wire  io_in_3_bits_exceptionVec_1;
  wire  io_in_3_bits_exceptionVec_2;
  wire  io_in_3_bits_exceptionVec_4;
  wire  io_in_3_bits_exceptionVec_5;
  wire  io_in_3_bits_exceptionVec_6;
  wire  io_in_3_bits_exceptionVec_7;
  wire  io_in_3_bits_exceptionVec_8;
  wire  io_in_3_bits_exceptionVec_9;
  wire  io_in_3_bits_exceptionVec_10;
  wire  io_in_3_bits_exceptionVec_11;
  wire  io_in_3_bits_exceptionVec_12;
  wire  io_in_3_bits_exceptionVec_13;
  wire  io_in_3_bits_exceptionVec_14;
  wire  io_in_3_bits_exceptionVec_15;
  wire  io_in_3_bits_exceptionVec_16;
  wire  io_in_3_bits_exceptionVec_17;
  wire  io_in_3_bits_exceptionVec_18;
  wire  io_in_3_bits_exceptionVec_19;
  wire  io_in_3_bits_exceptionVec_20;
  wire  io_in_3_bits_exceptionVec_21;
  wire  io_in_3_bits_exceptionVec_23;
  wire  io_in_3_bits_isFetchMalAddr;
  wire [3:0] io_in_3_bits_trigger;
  wire  io_in_3_bits_preDecodeInfo_isRVC;
  wire [1:0] io_in_3_bits_preDecodeInfo_brType;
  wire  io_in_3_bits_pred_taken;
  wire  io_in_3_bits_crossPageIPFFix;
  wire  io_in_3_bits_ftqPtr_flag;
  wire [5:0] io_in_3_bits_ftqPtr_value;
  wire [3:0] io_in_3_bits_ftqOffset;
  wire  io_in_3_bits_isLastInFtqEntry;
  wire  io_in_4_ready;
  wire  io_in_4_valid;
  wire [31:0] io_in_4_bits_instr;
  wire  io_in_4_bits_exceptionVec_0;
  wire  io_in_4_bits_exceptionVec_1;
  wire  io_in_4_bits_exceptionVec_2;
  wire  io_in_4_bits_exceptionVec_4;
  wire  io_in_4_bits_exceptionVec_5;
  wire  io_in_4_bits_exceptionVec_6;
  wire  io_in_4_bits_exceptionVec_7;
  wire  io_in_4_bits_exceptionVec_8;
  wire  io_in_4_bits_exceptionVec_9;
  wire  io_in_4_bits_exceptionVec_10;
  wire  io_in_4_bits_exceptionVec_11;
  wire  io_in_4_bits_exceptionVec_12;
  wire  io_in_4_bits_exceptionVec_13;
  wire  io_in_4_bits_exceptionVec_14;
  wire  io_in_4_bits_exceptionVec_15;
  wire  io_in_4_bits_exceptionVec_16;
  wire  io_in_4_bits_exceptionVec_17;
  wire  io_in_4_bits_exceptionVec_18;
  wire  io_in_4_bits_exceptionVec_19;
  wire  io_in_4_bits_exceptionVec_20;
  wire  io_in_4_bits_exceptionVec_21;
  wire  io_in_4_bits_exceptionVec_23;
  wire  io_in_4_bits_isFetchMalAddr;
  wire [3:0] io_in_4_bits_trigger;
  wire  io_in_4_bits_preDecodeInfo_isRVC;
  wire [1:0] io_in_4_bits_preDecodeInfo_brType;
  wire  io_in_4_bits_pred_taken;
  wire  io_in_4_bits_crossPageIPFFix;
  wire  io_in_4_bits_ftqPtr_flag;
  wire [5:0] io_in_4_bits_ftqPtr_value;
  wire [3:0] io_in_4_bits_ftqOffset;
  wire  io_in_4_bits_isLastInFtqEntry;
  wire  io_in_5_ready;
  wire  io_in_5_valid;
  wire [31:0] io_in_5_bits_instr;
  wire  io_in_5_bits_exceptionVec_0;
  wire  io_in_5_bits_exceptionVec_1;
  wire  io_in_5_bits_exceptionVec_2;
  wire  io_in_5_bits_exceptionVec_4;
  wire  io_in_5_bits_exceptionVec_5;
  wire  io_in_5_bits_exceptionVec_6;
  wire  io_in_5_bits_exceptionVec_7;
  wire  io_in_5_bits_exceptionVec_8;
  wire  io_in_5_bits_exceptionVec_9;
  wire  io_in_5_bits_exceptionVec_10;
  wire  io_in_5_bits_exceptionVec_11;
  wire  io_in_5_bits_exceptionVec_12;
  wire  io_in_5_bits_exceptionVec_13;
  wire  io_in_5_bits_exceptionVec_14;
  wire  io_in_5_bits_exceptionVec_15;
  wire  io_in_5_bits_exceptionVec_16;
  wire  io_in_5_bits_exceptionVec_17;
  wire  io_in_5_bits_exceptionVec_18;
  wire  io_in_5_bits_exceptionVec_19;
  wire  io_in_5_bits_exceptionVec_20;
  wire  io_in_5_bits_exceptionVec_21;
  wire  io_in_5_bits_exceptionVec_23;
  wire  io_in_5_bits_isFetchMalAddr;
  wire [3:0] io_in_5_bits_trigger;
  wire  io_in_5_bits_preDecodeInfo_isRVC;
  wire [1:0] io_in_5_bits_preDecodeInfo_brType;
  wire  io_in_5_bits_pred_taken;
  wire  io_in_5_bits_crossPageIPFFix;
  wire  io_in_5_bits_ftqPtr_flag;
  wire [5:0] io_in_5_bits_ftqPtr_value;
  wire [3:0] io_in_5_bits_ftqOffset;
  wire  io_in_5_bits_isLastInFtqEntry;
  wire  io_out_0_ready;
  wire  io_out_0_valid;
  wire [31:0] io_out_0_bits_instr;
  wire  io_out_0_bits_exceptionVec_0;
  wire  io_out_0_bits_exceptionVec_1;
  wire  io_out_0_bits_exceptionVec_2;
  wire  io_out_0_bits_exceptionVec_3;
  wire  io_out_0_bits_exceptionVec_4;
  wire  io_out_0_bits_exceptionVec_5;
  wire  io_out_0_bits_exceptionVec_6;
  wire  io_out_0_bits_exceptionVec_7;
  wire  io_out_0_bits_exceptionVec_8;
  wire  io_out_0_bits_exceptionVec_9;
  wire  io_out_0_bits_exceptionVec_10;
  wire  io_out_0_bits_exceptionVec_11;
  wire  io_out_0_bits_exceptionVec_12;
  wire  io_out_0_bits_exceptionVec_13;
  wire  io_out_0_bits_exceptionVec_14;
  wire  io_out_0_bits_exceptionVec_15;
  wire  io_out_0_bits_exceptionVec_16;
  wire  io_out_0_bits_exceptionVec_17;
  wire  io_out_0_bits_exceptionVec_18;
  wire  io_out_0_bits_exceptionVec_19;
  wire  io_out_0_bits_exceptionVec_20;
  wire  io_out_0_bits_exceptionVec_21;
  wire  io_out_0_bits_exceptionVec_22;
  wire  io_out_0_bits_exceptionVec_23;
  wire  io_out_0_bits_isFetchMalAddr;
  wire [3:0] io_out_0_bits_trigger;
  wire  io_out_0_bits_preDecodeInfo_isRVC;
  wire [1:0] io_out_0_bits_preDecodeInfo_brType;
  wire  io_out_0_bits_pred_taken;
  wire  io_out_0_bits_crossPageIPFFix;
  wire  io_out_0_bits_ftqPtr_flag;
  wire [5:0] io_out_0_bits_ftqPtr_value;
  wire [3:0] io_out_0_bits_ftqOffset;
  wire [3:0] io_out_0_bits_srcType_0;
  wire [3:0] io_out_0_bits_srcType_1;
  wire [3:0] io_out_0_bits_srcType_2;
  wire [3:0] io_out_0_bits_srcType_3;
  wire [3:0] io_out_0_bits_srcType_4;
  wire [5:0] io_out_0_bits_lsrc_0;
  wire [5:0] io_out_0_bits_lsrc_1;
  wire [5:0] io_out_0_bits_lsrc_2;
  wire [5:0] io_out_0_bits_ldest;
  wire [34:0] io_out_0_bits_fuType;
  wire [8:0] io_out_0_bits_fuOpType;
  wire  io_out_0_bits_rfWen;
  wire  io_out_0_bits_fpWen;
  wire  io_out_0_bits_vecWen;
  wire  io_out_0_bits_v0Wen;
  wire  io_out_0_bits_vlWen;
  wire  io_out_0_bits_isXSTrap;
  wire  io_out_0_bits_waitForward;
  wire  io_out_0_bits_blockBackward;
  wire  io_out_0_bits_flushPipe;
  wire  io_out_0_bits_canRobCompress;
  wire [3:0] io_out_0_bits_selImm;
  wire [21:0] io_out_0_bits_imm;
  wire [1:0] io_out_0_bits_fpu_typeTagOut;
  wire  io_out_0_bits_fpu_wflags;
  wire [1:0] io_out_0_bits_fpu_typ;
  wire [1:0] io_out_0_bits_fpu_fmt;
  wire [2:0] io_out_0_bits_fpu_rm;
  wire  io_out_0_bits_vpu_vill;
  wire  io_out_0_bits_vpu_vma;
  wire  io_out_0_bits_vpu_vta;
  wire [1:0] io_out_0_bits_vpu_vsew;
  wire [2:0] io_out_0_bits_vpu_vlmul;
  wire  io_out_0_bits_vpu_specVill;
  wire  io_out_0_bits_vpu_specVma;
  wire  io_out_0_bits_vpu_specVta;
  wire [1:0] io_out_0_bits_vpu_specVsew;
  wire [2:0] io_out_0_bits_vpu_specVlmul;
  wire  io_out_0_bits_vpu_vm;
  wire [7:0] io_out_0_bits_vpu_vstart;
  wire  io_out_0_bits_vpu_fpu_isFoldTo1_2;
  wire  io_out_0_bits_vpu_fpu_isFoldTo1_4;
  wire  io_out_0_bits_vpu_fpu_isFoldTo1_8;
  wire [2:0] io_out_0_bits_vpu_nf;
  wire [1:0] io_out_0_bits_vpu_veew;
  wire  io_out_0_bits_vpu_isExt;
  wire  io_out_0_bits_vpu_isNarrow;
  wire  io_out_0_bits_vpu_isDstMask;
  wire  io_out_0_bits_vpu_isOpMask;
  wire  io_out_0_bits_vpu_isDependOldVd;
  wire  io_out_0_bits_vpu_isWritePartVd;
  wire  io_out_0_bits_vpu_isVleff;
  wire  io_out_0_bits_vlsInstr;
  wire  io_out_0_bits_wfflags;
  wire  io_out_0_bits_isMove;
  wire [6:0] io_out_0_bits_uopIdx;
  wire [5:0] io_out_0_bits_uopSplitType;
  wire  io_out_0_bits_isVset;
  wire  io_out_0_bits_firstUop;
  wire  io_out_0_bits_lastUop;
  wire [6:0] io_out_0_bits_numWB;
  wire [2:0] io_out_0_bits_commitType;
  wire  io_out_1_ready;
  wire  io_out_1_valid;
  wire [31:0] io_out_1_bits_instr;
  wire  io_out_1_bits_exceptionVec_0;
  wire  io_out_1_bits_exceptionVec_1;
  wire  io_out_1_bits_exceptionVec_2;
  wire  io_out_1_bits_exceptionVec_3;
  wire  io_out_1_bits_exceptionVec_4;
  wire  io_out_1_bits_exceptionVec_5;
  wire  io_out_1_bits_exceptionVec_6;
  wire  io_out_1_bits_exceptionVec_7;
  wire  io_out_1_bits_exceptionVec_8;
  wire  io_out_1_bits_exceptionVec_9;
  wire  io_out_1_bits_exceptionVec_10;
  wire  io_out_1_bits_exceptionVec_11;
  wire  io_out_1_bits_exceptionVec_12;
  wire  io_out_1_bits_exceptionVec_13;
  wire  io_out_1_bits_exceptionVec_14;
  wire  io_out_1_bits_exceptionVec_15;
  wire  io_out_1_bits_exceptionVec_16;
  wire  io_out_1_bits_exceptionVec_17;
  wire  io_out_1_bits_exceptionVec_18;
  wire  io_out_1_bits_exceptionVec_19;
  wire  io_out_1_bits_exceptionVec_20;
  wire  io_out_1_bits_exceptionVec_21;
  wire  io_out_1_bits_exceptionVec_22;
  wire  io_out_1_bits_exceptionVec_23;
  wire  io_out_1_bits_isFetchMalAddr;
  wire [3:0] io_out_1_bits_trigger;
  wire  io_out_1_bits_preDecodeInfo_isRVC;
  wire [1:0] io_out_1_bits_preDecodeInfo_brType;
  wire  io_out_1_bits_pred_taken;
  wire  io_out_1_bits_crossPageIPFFix;
  wire  io_out_1_bits_ftqPtr_flag;
  wire [5:0] io_out_1_bits_ftqPtr_value;
  wire [3:0] io_out_1_bits_ftqOffset;
  wire [3:0] io_out_1_bits_srcType_0;
  wire [3:0] io_out_1_bits_srcType_1;
  wire [3:0] io_out_1_bits_srcType_2;
  wire [3:0] io_out_1_bits_srcType_3;
  wire [3:0] io_out_1_bits_srcType_4;
  wire [5:0] io_out_1_bits_lsrc_0;
  wire [5:0] io_out_1_bits_lsrc_1;
  wire [5:0] io_out_1_bits_lsrc_2;
  wire [5:0] io_out_1_bits_ldest;
  wire [34:0] io_out_1_bits_fuType;
  wire [8:0] io_out_1_bits_fuOpType;
  wire  io_out_1_bits_rfWen;
  wire  io_out_1_bits_fpWen;
  wire  io_out_1_bits_vecWen;
  wire  io_out_1_bits_v0Wen;
  wire  io_out_1_bits_vlWen;
  wire  io_out_1_bits_isXSTrap;
  wire  io_out_1_bits_waitForward;
  wire  io_out_1_bits_blockBackward;
  wire  io_out_1_bits_flushPipe;
  wire  io_out_1_bits_canRobCompress;
  wire [3:0] io_out_1_bits_selImm;
  wire [21:0] io_out_1_bits_imm;
  wire [1:0] io_out_1_bits_fpu_typeTagOut;
  wire  io_out_1_bits_fpu_wflags;
  wire [1:0] io_out_1_bits_fpu_typ;
  wire [1:0] io_out_1_bits_fpu_fmt;
  wire [2:0] io_out_1_bits_fpu_rm;
  wire  io_out_1_bits_vpu_vill;
  wire  io_out_1_bits_vpu_vma;
  wire  io_out_1_bits_vpu_vta;
  wire [1:0] io_out_1_bits_vpu_vsew;
  wire [2:0] io_out_1_bits_vpu_vlmul;
  wire  io_out_1_bits_vpu_specVill;
  wire  io_out_1_bits_vpu_specVma;
  wire  io_out_1_bits_vpu_specVta;
  wire [1:0] io_out_1_bits_vpu_specVsew;
  wire [2:0] io_out_1_bits_vpu_specVlmul;
  wire  io_out_1_bits_vpu_vm;
  wire [7:0] io_out_1_bits_vpu_vstart;
  wire  io_out_1_bits_vpu_fpu_isFoldTo1_2;
  wire  io_out_1_bits_vpu_fpu_isFoldTo1_4;
  wire  io_out_1_bits_vpu_fpu_isFoldTo1_8;
  wire [2:0] io_out_1_bits_vpu_nf;
  wire [1:0] io_out_1_bits_vpu_veew;
  wire  io_out_1_bits_vpu_isExt;
  wire  io_out_1_bits_vpu_isNarrow;
  wire  io_out_1_bits_vpu_isDstMask;
  wire  io_out_1_bits_vpu_isOpMask;
  wire  io_out_1_bits_vpu_isDependOldVd;
  wire  io_out_1_bits_vpu_isWritePartVd;
  wire  io_out_1_bits_vpu_isVleff;
  wire  io_out_1_bits_vlsInstr;
  wire  io_out_1_bits_wfflags;
  wire  io_out_1_bits_isMove;
  wire [6:0] io_out_1_bits_uopIdx;
  wire [5:0] io_out_1_bits_uopSplitType;
  wire  io_out_1_bits_isVset;
  wire  io_out_1_bits_firstUop;
  wire  io_out_1_bits_lastUop;
  wire [6:0] io_out_1_bits_numWB;
  wire [2:0] io_out_1_bits_commitType;
  wire  io_out_2_ready;
  wire  io_out_2_valid;
  wire [31:0] io_out_2_bits_instr;
  wire  io_out_2_bits_exceptionVec_0;
  wire  io_out_2_bits_exceptionVec_1;
  wire  io_out_2_bits_exceptionVec_2;
  wire  io_out_2_bits_exceptionVec_3;
  wire  io_out_2_bits_exceptionVec_4;
  wire  io_out_2_bits_exceptionVec_5;
  wire  io_out_2_bits_exceptionVec_6;
  wire  io_out_2_bits_exceptionVec_7;
  wire  io_out_2_bits_exceptionVec_8;
  wire  io_out_2_bits_exceptionVec_9;
  wire  io_out_2_bits_exceptionVec_10;
  wire  io_out_2_bits_exceptionVec_11;
  wire  io_out_2_bits_exceptionVec_12;
  wire  io_out_2_bits_exceptionVec_13;
  wire  io_out_2_bits_exceptionVec_14;
  wire  io_out_2_bits_exceptionVec_15;
  wire  io_out_2_bits_exceptionVec_16;
  wire  io_out_2_bits_exceptionVec_17;
  wire  io_out_2_bits_exceptionVec_18;
  wire  io_out_2_bits_exceptionVec_19;
  wire  io_out_2_bits_exceptionVec_20;
  wire  io_out_2_bits_exceptionVec_21;
  wire  io_out_2_bits_exceptionVec_22;
  wire  io_out_2_bits_exceptionVec_23;
  wire  io_out_2_bits_isFetchMalAddr;
  wire [3:0] io_out_2_bits_trigger;
  wire  io_out_2_bits_preDecodeInfo_isRVC;
  wire [1:0] io_out_2_bits_preDecodeInfo_brType;
  wire  io_out_2_bits_pred_taken;
  wire  io_out_2_bits_crossPageIPFFix;
  wire  io_out_2_bits_ftqPtr_flag;
  wire [5:0] io_out_2_bits_ftqPtr_value;
  wire [3:0] io_out_2_bits_ftqOffset;
  wire [3:0] io_out_2_bits_srcType_0;
  wire [3:0] io_out_2_bits_srcType_1;
  wire [3:0] io_out_2_bits_srcType_2;
  wire [3:0] io_out_2_bits_srcType_3;
  wire [3:0] io_out_2_bits_srcType_4;
  wire [5:0] io_out_2_bits_lsrc_0;
  wire [5:0] io_out_2_bits_lsrc_1;
  wire [5:0] io_out_2_bits_lsrc_2;
  wire [5:0] io_out_2_bits_ldest;
  wire [34:0] io_out_2_bits_fuType;
  wire [8:0] io_out_2_bits_fuOpType;
  wire  io_out_2_bits_rfWen;
  wire  io_out_2_bits_fpWen;
  wire  io_out_2_bits_vecWen;
  wire  io_out_2_bits_v0Wen;
  wire  io_out_2_bits_vlWen;
  wire  io_out_2_bits_isXSTrap;
  wire  io_out_2_bits_waitForward;
  wire  io_out_2_bits_blockBackward;
  wire  io_out_2_bits_flushPipe;
  wire  io_out_2_bits_canRobCompress;
  wire [3:0] io_out_2_bits_selImm;
  wire [21:0] io_out_2_bits_imm;
  wire [1:0] io_out_2_bits_fpu_typeTagOut;
  wire  io_out_2_bits_fpu_wflags;
  wire [1:0] io_out_2_bits_fpu_typ;
  wire [1:0] io_out_2_bits_fpu_fmt;
  wire [2:0] io_out_2_bits_fpu_rm;
  wire  io_out_2_bits_vpu_vill;
  wire  io_out_2_bits_vpu_vma;
  wire  io_out_2_bits_vpu_vta;
  wire [1:0] io_out_2_bits_vpu_vsew;
  wire [2:0] io_out_2_bits_vpu_vlmul;
  wire  io_out_2_bits_vpu_specVill;
  wire  io_out_2_bits_vpu_specVma;
  wire  io_out_2_bits_vpu_specVta;
  wire [1:0] io_out_2_bits_vpu_specVsew;
  wire [2:0] io_out_2_bits_vpu_specVlmul;
  wire  io_out_2_bits_vpu_vm;
  wire [7:0] io_out_2_bits_vpu_vstart;
  wire  io_out_2_bits_vpu_fpu_isFoldTo1_2;
  wire  io_out_2_bits_vpu_fpu_isFoldTo1_4;
  wire  io_out_2_bits_vpu_fpu_isFoldTo1_8;
  wire [2:0] io_out_2_bits_vpu_nf;
  wire [1:0] io_out_2_bits_vpu_veew;
  wire  io_out_2_bits_vpu_isExt;
  wire  io_out_2_bits_vpu_isNarrow;
  wire  io_out_2_bits_vpu_isDstMask;
  wire  io_out_2_bits_vpu_isOpMask;
  wire  io_out_2_bits_vpu_isDependOldVd;
  wire  io_out_2_bits_vpu_isWritePartVd;
  wire  io_out_2_bits_vpu_isVleff;
  wire  io_out_2_bits_vlsInstr;
  wire  io_out_2_bits_wfflags;
  wire  io_out_2_bits_isMove;
  wire [6:0] io_out_2_bits_uopIdx;
  wire [5:0] io_out_2_bits_uopSplitType;
  wire  io_out_2_bits_isVset;
  wire  io_out_2_bits_firstUop;
  wire  io_out_2_bits_lastUop;
  wire [6:0] io_out_2_bits_numWB;
  wire [2:0] io_out_2_bits_commitType;
  wire  io_out_3_ready;
  wire  io_out_3_valid;
  wire [31:0] io_out_3_bits_instr;
  wire  io_out_3_bits_exceptionVec_0;
  wire  io_out_3_bits_exceptionVec_1;
  wire  io_out_3_bits_exceptionVec_2;
  wire  io_out_3_bits_exceptionVec_3;
  wire  io_out_3_bits_exceptionVec_4;
  wire  io_out_3_bits_exceptionVec_5;
  wire  io_out_3_bits_exceptionVec_6;
  wire  io_out_3_bits_exceptionVec_7;
  wire  io_out_3_bits_exceptionVec_8;
  wire  io_out_3_bits_exceptionVec_9;
  wire  io_out_3_bits_exceptionVec_10;
  wire  io_out_3_bits_exceptionVec_11;
  wire  io_out_3_bits_exceptionVec_12;
  wire  io_out_3_bits_exceptionVec_13;
  wire  io_out_3_bits_exceptionVec_14;
  wire  io_out_3_bits_exceptionVec_15;
  wire  io_out_3_bits_exceptionVec_16;
  wire  io_out_3_bits_exceptionVec_17;
  wire  io_out_3_bits_exceptionVec_18;
  wire  io_out_3_bits_exceptionVec_19;
  wire  io_out_3_bits_exceptionVec_20;
  wire  io_out_3_bits_exceptionVec_21;
  wire  io_out_3_bits_exceptionVec_22;
  wire  io_out_3_bits_exceptionVec_23;
  wire  io_out_3_bits_isFetchMalAddr;
  wire [3:0] io_out_3_bits_trigger;
  wire  io_out_3_bits_preDecodeInfo_isRVC;
  wire [1:0] io_out_3_bits_preDecodeInfo_brType;
  wire  io_out_3_bits_pred_taken;
  wire  io_out_3_bits_crossPageIPFFix;
  wire  io_out_3_bits_ftqPtr_flag;
  wire [5:0] io_out_3_bits_ftqPtr_value;
  wire [3:0] io_out_3_bits_ftqOffset;
  wire [3:0] io_out_3_bits_srcType_0;
  wire [3:0] io_out_3_bits_srcType_1;
  wire [3:0] io_out_3_bits_srcType_2;
  wire [3:0] io_out_3_bits_srcType_3;
  wire [3:0] io_out_3_bits_srcType_4;
  wire [5:0] io_out_3_bits_lsrc_0;
  wire [5:0] io_out_3_bits_lsrc_1;
  wire [5:0] io_out_3_bits_lsrc_2;
  wire [5:0] io_out_3_bits_ldest;
  wire [34:0] io_out_3_bits_fuType;
  wire [8:0] io_out_3_bits_fuOpType;
  wire  io_out_3_bits_rfWen;
  wire  io_out_3_bits_fpWen;
  wire  io_out_3_bits_vecWen;
  wire  io_out_3_bits_v0Wen;
  wire  io_out_3_bits_vlWen;
  wire  io_out_3_bits_isXSTrap;
  wire  io_out_3_bits_waitForward;
  wire  io_out_3_bits_blockBackward;
  wire  io_out_3_bits_flushPipe;
  wire  io_out_3_bits_canRobCompress;
  wire [3:0] io_out_3_bits_selImm;
  wire [21:0] io_out_3_bits_imm;
  wire [1:0] io_out_3_bits_fpu_typeTagOut;
  wire  io_out_3_bits_fpu_wflags;
  wire [1:0] io_out_3_bits_fpu_typ;
  wire [1:0] io_out_3_bits_fpu_fmt;
  wire [2:0] io_out_3_bits_fpu_rm;
  wire  io_out_3_bits_vpu_vill;
  wire  io_out_3_bits_vpu_vma;
  wire  io_out_3_bits_vpu_vta;
  wire [1:0] io_out_3_bits_vpu_vsew;
  wire [2:0] io_out_3_bits_vpu_vlmul;
  wire  io_out_3_bits_vpu_specVill;
  wire  io_out_3_bits_vpu_specVma;
  wire  io_out_3_bits_vpu_specVta;
  wire [1:0] io_out_3_bits_vpu_specVsew;
  wire [2:0] io_out_3_bits_vpu_specVlmul;
  wire  io_out_3_bits_vpu_vm;
  wire [7:0] io_out_3_bits_vpu_vstart;
  wire  io_out_3_bits_vpu_fpu_isFoldTo1_2;
  wire  io_out_3_bits_vpu_fpu_isFoldTo1_4;
  wire  io_out_3_bits_vpu_fpu_isFoldTo1_8;
  wire [2:0] io_out_3_bits_vpu_nf;
  wire [1:0] io_out_3_bits_vpu_veew;
  wire  io_out_3_bits_vpu_isExt;
  wire  io_out_3_bits_vpu_isNarrow;
  wire  io_out_3_bits_vpu_isDstMask;
  wire  io_out_3_bits_vpu_isOpMask;
  wire  io_out_3_bits_vpu_isDependOldVd;
  wire  io_out_3_bits_vpu_isWritePartVd;
  wire  io_out_3_bits_vpu_isVleff;
  wire  io_out_3_bits_vlsInstr;
  wire  io_out_3_bits_wfflags;
  wire  io_out_3_bits_isMove;
  wire [6:0] io_out_3_bits_uopIdx;
  wire [5:0] io_out_3_bits_uopSplitType;
  wire  io_out_3_bits_isVset;
  wire  io_out_3_bits_firstUop;
  wire  io_out_3_bits_lastUop;
  wire [6:0] io_out_3_bits_numWB;
  wire [2:0] io_out_3_bits_commitType;
  wire  io_out_4_ready;
  wire  io_out_4_valid;
  wire [31:0] io_out_4_bits_instr;
  wire  io_out_4_bits_exceptionVec_0;
  wire  io_out_4_bits_exceptionVec_1;
  wire  io_out_4_bits_exceptionVec_2;
  wire  io_out_4_bits_exceptionVec_3;
  wire  io_out_4_bits_exceptionVec_4;
  wire  io_out_4_bits_exceptionVec_5;
  wire  io_out_4_bits_exceptionVec_6;
  wire  io_out_4_bits_exceptionVec_7;
  wire  io_out_4_bits_exceptionVec_8;
  wire  io_out_4_bits_exceptionVec_9;
  wire  io_out_4_bits_exceptionVec_10;
  wire  io_out_4_bits_exceptionVec_11;
  wire  io_out_4_bits_exceptionVec_12;
  wire  io_out_4_bits_exceptionVec_13;
  wire  io_out_4_bits_exceptionVec_14;
  wire  io_out_4_bits_exceptionVec_15;
  wire  io_out_4_bits_exceptionVec_16;
  wire  io_out_4_bits_exceptionVec_17;
  wire  io_out_4_bits_exceptionVec_18;
  wire  io_out_4_bits_exceptionVec_19;
  wire  io_out_4_bits_exceptionVec_20;
  wire  io_out_4_bits_exceptionVec_21;
  wire  io_out_4_bits_exceptionVec_22;
  wire  io_out_4_bits_exceptionVec_23;
  wire  io_out_4_bits_isFetchMalAddr;
  wire [3:0] io_out_4_bits_trigger;
  wire  io_out_4_bits_preDecodeInfo_isRVC;
  wire [1:0] io_out_4_bits_preDecodeInfo_brType;
  wire  io_out_4_bits_pred_taken;
  wire  io_out_4_bits_crossPageIPFFix;
  wire  io_out_4_bits_ftqPtr_flag;
  wire [5:0] io_out_4_bits_ftqPtr_value;
  wire [3:0] io_out_4_bits_ftqOffset;
  wire [3:0] io_out_4_bits_srcType_0;
  wire [3:0] io_out_4_bits_srcType_1;
  wire [3:0] io_out_4_bits_srcType_2;
  wire [3:0] io_out_4_bits_srcType_3;
  wire [3:0] io_out_4_bits_srcType_4;
  wire [5:0] io_out_4_bits_lsrc_0;
  wire [5:0] io_out_4_bits_lsrc_1;
  wire [5:0] io_out_4_bits_lsrc_2;
  wire [5:0] io_out_4_bits_ldest;
  wire [34:0] io_out_4_bits_fuType;
  wire [8:0] io_out_4_bits_fuOpType;
  wire  io_out_4_bits_rfWen;
  wire  io_out_4_bits_fpWen;
  wire  io_out_4_bits_vecWen;
  wire  io_out_4_bits_v0Wen;
  wire  io_out_4_bits_vlWen;
  wire  io_out_4_bits_isXSTrap;
  wire  io_out_4_bits_waitForward;
  wire  io_out_4_bits_blockBackward;
  wire  io_out_4_bits_flushPipe;
  wire  io_out_4_bits_canRobCompress;
  wire [3:0] io_out_4_bits_selImm;
  wire [21:0] io_out_4_bits_imm;
  wire [1:0] io_out_4_bits_fpu_typeTagOut;
  wire  io_out_4_bits_fpu_wflags;
  wire [1:0] io_out_4_bits_fpu_typ;
  wire [1:0] io_out_4_bits_fpu_fmt;
  wire [2:0] io_out_4_bits_fpu_rm;
  wire  io_out_4_bits_vpu_vill;
  wire  io_out_4_bits_vpu_vma;
  wire  io_out_4_bits_vpu_vta;
  wire [1:0] io_out_4_bits_vpu_vsew;
  wire [2:0] io_out_4_bits_vpu_vlmul;
  wire  io_out_4_bits_vpu_specVill;
  wire  io_out_4_bits_vpu_specVma;
  wire  io_out_4_bits_vpu_specVta;
  wire [1:0] io_out_4_bits_vpu_specVsew;
  wire [2:0] io_out_4_bits_vpu_specVlmul;
  wire  io_out_4_bits_vpu_vm;
  wire [7:0] io_out_4_bits_vpu_vstart;
  wire  io_out_4_bits_vpu_fpu_isFoldTo1_2;
  wire  io_out_4_bits_vpu_fpu_isFoldTo1_4;
  wire  io_out_4_bits_vpu_fpu_isFoldTo1_8;
  wire [2:0] io_out_4_bits_vpu_nf;
  wire [1:0] io_out_4_bits_vpu_veew;
  wire  io_out_4_bits_vpu_isExt;
  wire  io_out_4_bits_vpu_isNarrow;
  wire  io_out_4_bits_vpu_isDstMask;
  wire  io_out_4_bits_vpu_isOpMask;
  wire  io_out_4_bits_vpu_isDependOldVd;
  wire  io_out_4_bits_vpu_isWritePartVd;
  wire  io_out_4_bits_vpu_isVleff;
  wire  io_out_4_bits_vlsInstr;
  wire  io_out_4_bits_wfflags;
  wire  io_out_4_bits_isMove;
  wire [6:0] io_out_4_bits_uopIdx;
  wire [5:0] io_out_4_bits_uopSplitType;
  wire  io_out_4_bits_isVset;
  wire  io_out_4_bits_firstUop;
  wire  io_out_4_bits_lastUop;
  wire [6:0] io_out_4_bits_numWB;
  wire [2:0] io_out_4_bits_commitType;
  wire  io_out_5_ready;
  wire  io_out_5_valid;
  wire [31:0] io_out_5_bits_instr;
  wire  io_out_5_bits_exceptionVec_0;
  wire  io_out_5_bits_exceptionVec_1;
  wire  io_out_5_bits_exceptionVec_2;
  wire  io_out_5_bits_exceptionVec_3;
  wire  io_out_5_bits_exceptionVec_4;
  wire  io_out_5_bits_exceptionVec_5;
  wire  io_out_5_bits_exceptionVec_6;
  wire  io_out_5_bits_exceptionVec_7;
  wire  io_out_5_bits_exceptionVec_8;
  wire  io_out_5_bits_exceptionVec_9;
  wire  io_out_5_bits_exceptionVec_10;
  wire  io_out_5_bits_exceptionVec_11;
  wire  io_out_5_bits_exceptionVec_12;
  wire  io_out_5_bits_exceptionVec_13;
  wire  io_out_5_bits_exceptionVec_14;
  wire  io_out_5_bits_exceptionVec_15;
  wire  io_out_5_bits_exceptionVec_16;
  wire  io_out_5_bits_exceptionVec_17;
  wire  io_out_5_bits_exceptionVec_18;
  wire  io_out_5_bits_exceptionVec_19;
  wire  io_out_5_bits_exceptionVec_20;
  wire  io_out_5_bits_exceptionVec_21;
  wire  io_out_5_bits_exceptionVec_22;
  wire  io_out_5_bits_exceptionVec_23;
  wire  io_out_5_bits_isFetchMalAddr;
  wire [3:0] io_out_5_bits_trigger;
  wire  io_out_5_bits_preDecodeInfo_isRVC;
  wire [1:0] io_out_5_bits_preDecodeInfo_brType;
  wire  io_out_5_bits_pred_taken;
  wire  io_out_5_bits_crossPageIPFFix;
  wire  io_out_5_bits_ftqPtr_flag;
  wire [5:0] io_out_5_bits_ftqPtr_value;
  wire [3:0] io_out_5_bits_ftqOffset;
  wire [3:0] io_out_5_bits_srcType_0;
  wire [3:0] io_out_5_bits_srcType_1;
  wire [3:0] io_out_5_bits_srcType_2;
  wire [3:0] io_out_5_bits_srcType_3;
  wire [3:0] io_out_5_bits_srcType_4;
  wire [5:0] io_out_5_bits_lsrc_0;
  wire [5:0] io_out_5_bits_lsrc_1;
  wire [5:0] io_out_5_bits_lsrc_2;
  wire [5:0] io_out_5_bits_ldest;
  wire [34:0] io_out_5_bits_fuType;
  wire [8:0] io_out_5_bits_fuOpType;
  wire  io_out_5_bits_rfWen;
  wire  io_out_5_bits_fpWen;
  wire  io_out_5_bits_vecWen;
  wire  io_out_5_bits_v0Wen;
  wire  io_out_5_bits_vlWen;
  wire  io_out_5_bits_isXSTrap;
  wire  io_out_5_bits_waitForward;
  wire  io_out_5_bits_blockBackward;
  wire  io_out_5_bits_flushPipe;
  wire  io_out_5_bits_canRobCompress;
  wire [3:0] io_out_5_bits_selImm;
  wire [21:0] io_out_5_bits_imm;
  wire [1:0] io_out_5_bits_fpu_typeTagOut;
  wire  io_out_5_bits_fpu_wflags;
  wire [1:0] io_out_5_bits_fpu_typ;
  wire [1:0] io_out_5_bits_fpu_fmt;
  wire [2:0] io_out_5_bits_fpu_rm;
  wire  io_out_5_bits_vpu_vill;
  wire  io_out_5_bits_vpu_vma;
  wire  io_out_5_bits_vpu_vta;
  wire [1:0] io_out_5_bits_vpu_vsew;
  wire [2:0] io_out_5_bits_vpu_vlmul;
  wire  io_out_5_bits_vpu_specVill;
  wire  io_out_5_bits_vpu_specVma;
  wire  io_out_5_bits_vpu_specVta;
  wire [1:0] io_out_5_bits_vpu_specVsew;
  wire [2:0] io_out_5_bits_vpu_specVlmul;
  wire  io_out_5_bits_vpu_vm;
  wire [7:0] io_out_5_bits_vpu_vstart;
  wire  io_out_5_bits_vpu_fpu_isFoldTo1_2;
  wire  io_out_5_bits_vpu_fpu_isFoldTo1_4;
  wire  io_out_5_bits_vpu_fpu_isFoldTo1_8;
  wire [2:0] io_out_5_bits_vpu_nf;
  wire [1:0] io_out_5_bits_vpu_veew;
  wire  io_out_5_bits_vpu_isExt;
  wire  io_out_5_bits_vpu_isNarrow;
  wire  io_out_5_bits_vpu_isDstMask;
  wire  io_out_5_bits_vpu_isOpMask;
  wire  io_out_5_bits_vpu_isDependOldVd;
  wire  io_out_5_bits_vpu_isWritePartVd;
  wire  io_out_5_bits_vpu_isVleff;
  wire  io_out_5_bits_vlsInstr;
  wire  io_out_5_bits_wfflags;
  wire  io_out_5_bits_isMove;
  wire [6:0] io_out_5_bits_uopIdx;
  wire [5:0] io_out_5_bits_uopSplitType;
  wire  io_out_5_bits_isVset;
  wire  io_out_5_bits_firstUop;
  wire  io_out_5_bits_lastUop;
  wire [6:0] io_out_5_bits_numWB;
  wire [2:0] io_out_5_bits_commitType;
  wire  io_intRat_0_0_hold;
  wire [31:0] io_intRat_0_0_addr;
  wire  io_intRat_0_1_hold;
  wire [31:0] io_intRat_0_1_addr;
  wire  io_intRat_1_0_hold;
  wire [31:0] io_intRat_1_0_addr;
  wire  io_intRat_1_1_hold;
  wire [31:0] io_intRat_1_1_addr;
  wire  io_intRat_2_0_hold;
  wire [31:0] io_intRat_2_0_addr;
  wire  io_intRat_2_1_hold;
  wire [31:0] io_intRat_2_1_addr;
  wire  io_intRat_3_0_hold;
  wire [31:0] io_intRat_3_0_addr;
  wire  io_intRat_3_1_hold;
  wire [31:0] io_intRat_3_1_addr;
  wire  io_intRat_4_0_hold;
  wire [31:0] io_intRat_4_0_addr;
  wire  io_intRat_4_1_hold;
  wire [31:0] io_intRat_4_1_addr;
  wire  io_intRat_5_0_hold;
  wire [31:0] io_intRat_5_0_addr;
  wire  io_intRat_5_1_hold;
  wire [31:0] io_intRat_5_1_addr;
  wire  io_fpRat_0_0_hold;
  wire [33:0] io_fpRat_0_0_addr;
  wire  io_fpRat_0_1_hold;
  wire [33:0] io_fpRat_0_1_addr;
  wire  io_fpRat_0_2_hold;
  wire [33:0] io_fpRat_0_2_addr;
  wire  io_fpRat_1_0_hold;
  wire [33:0] io_fpRat_1_0_addr;
  wire  io_fpRat_1_1_hold;
  wire [33:0] io_fpRat_1_1_addr;
  wire  io_fpRat_1_2_hold;
  wire [33:0] io_fpRat_1_2_addr;
  wire  io_fpRat_2_0_hold;
  wire [33:0] io_fpRat_2_0_addr;
  wire  io_fpRat_2_1_hold;
  wire [33:0] io_fpRat_2_1_addr;
  wire  io_fpRat_2_2_hold;
  wire [33:0] io_fpRat_2_2_addr;
  wire  io_fpRat_3_0_hold;
  wire [33:0] io_fpRat_3_0_addr;
  wire  io_fpRat_3_1_hold;
  wire [33:0] io_fpRat_3_1_addr;
  wire  io_fpRat_3_2_hold;
  wire [33:0] io_fpRat_3_2_addr;
  wire  io_fpRat_4_0_hold;
  wire [33:0] io_fpRat_4_0_addr;
  wire  io_fpRat_4_1_hold;
  wire [33:0] io_fpRat_4_1_addr;
  wire  io_fpRat_4_2_hold;
  wire [33:0] io_fpRat_4_2_addr;
  wire  io_fpRat_5_0_hold;
  wire [33:0] io_fpRat_5_0_addr;
  wire  io_fpRat_5_1_hold;
  wire [33:0] io_fpRat_5_1_addr;
  wire  io_fpRat_5_2_hold;
  wire [33:0] io_fpRat_5_2_addr;
  wire  io_vecRat_0_0_hold;
  wire [46:0] io_vecRat_0_0_addr;
  wire  io_vecRat_0_1_hold;
  wire [46:0] io_vecRat_0_1_addr;
  wire  io_vecRat_0_2_hold;
  wire [46:0] io_vecRat_0_2_addr;
  wire  io_vecRat_1_0_hold;
  wire [46:0] io_vecRat_1_0_addr;
  wire  io_vecRat_1_1_hold;
  wire [46:0] io_vecRat_1_1_addr;
  wire  io_vecRat_1_2_hold;
  wire [46:0] io_vecRat_1_2_addr;
  wire  io_vecRat_2_0_hold;
  wire [46:0] io_vecRat_2_0_addr;
  wire  io_vecRat_2_1_hold;
  wire [46:0] io_vecRat_2_1_addr;
  wire  io_vecRat_2_2_hold;
  wire [46:0] io_vecRat_2_2_addr;
  wire  io_vecRat_3_0_hold;
  wire [46:0] io_vecRat_3_0_addr;
  wire  io_vecRat_3_1_hold;
  wire [46:0] io_vecRat_3_1_addr;
  wire  io_vecRat_3_2_hold;
  wire [46:0] io_vecRat_3_2_addr;
  wire  io_vecRat_4_0_hold;
  wire [46:0] io_vecRat_4_0_addr;
  wire  io_vecRat_4_1_hold;
  wire [46:0] io_vecRat_4_1_addr;
  wire  io_vecRat_4_2_hold;
  wire [46:0] io_vecRat_4_2_addr;
  wire  io_vecRat_5_0_hold;
  wire [46:0] io_vecRat_5_0_addr;
  wire  io_vecRat_5_1_hold;
  wire [46:0] io_vecRat_5_1_addr;
  wire  io_vecRat_5_2_hold;
  wire [46:0] io_vecRat_5_2_addr;
  wire  io_csrCtrl_singlestep;
  wire  io_fromCSR_illegalInst_sfenceVMA;
  wire  io_fromCSR_illegalInst_sfencePart;
  wire  io_fromCSR_illegalInst_hfenceGVMA;
  wire  io_fromCSR_illegalInst_hfenceVVMA;
  wire  io_fromCSR_illegalInst_hlsv;
  wire  io_fromCSR_illegalInst_fsIsOff;
  wire  io_fromCSR_illegalInst_vsIsOff;
  wire  io_fromCSR_illegalInst_wfi;
  wire  io_fromCSR_illegalInst_frm;
  wire  io_fromCSR_illegalInst_cboZ;
  wire  io_fromCSR_illegalInst_cboCF;
  wire  io_fromCSR_illegalInst_cboI;
  wire  io_fromCSR_virtualInst_sfenceVMA;
  wire  io_fromCSR_virtualInst_sfencePart;
  wire  io_fromCSR_virtualInst_hfence;
  wire  io_fromCSR_virtualInst_hlsv;
  wire  io_fromCSR_virtualInst_wfi;
  wire  io_fromCSR_virtualInst_cboZ;
  wire  io_fromCSR_virtualInst_cboCF;
  wire  io_fromCSR_virtualInst_cboI;
  wire  io_fromCSR_special_cboI2F;
  wire  io_fusion_0;
  wire  io_fusion_1;
  wire  io_fusion_2;
  wire  io_fusion_3;
  wire  io_fusion_4;
  wire  io_fromRob_isResumeVType;
  wire  io_fromRob_walkToArchVType;
  wire  io_fromRob_commitVType_vtype_valid;
  wire  io_fromRob_commitVType_vtype_bits_illegal;
  wire  io_fromRob_commitVType_vtype_bits_vma;
  wire  io_fromRob_commitVType_vtype_bits_vta;
  wire [1:0] io_fromRob_commitVType_vtype_bits_vsew;
  wire [2:0] io_fromRob_commitVType_vtype_bits_vlmul;
  wire  io_fromRob_commitVType_hasVsetvl;
  wire  io_fromRob_walkVType_valid;
  wire  io_fromRob_walkVType_bits_illegal;
  wire  io_fromRob_walkVType_bits_vma;
  wire  io_fromRob_walkVType_bits_vta;
  wire [1:0] io_fromRob_walkVType_bits_vsew;
  wire [2:0] io_fromRob_walkVType_bits_vlmul;
  wire  io_vsetvlVType_illegal;
  wire  io_vsetvlVType_vma;
  wire  io_vsetvlVType_vta;
  wire [1:0] io_vsetvlVType_vsew;
  wire [2:0] io_vsetvlVType_vlmul;
  wire [7:0] io_vstart;
  wire  io_toCSR_trapInstInfo_valid;
  wire [31:0] io_toCSR_trapInstInfo_bits_instr;
  wire  io_toCSR_trapInstInfo_bits_ftqPtr_flag;
  wire [5:0] io_toCSR_trapInstInfo_bits_ftqPtr_value;
  wire [3:0] io_toCSR_trapInstInfo_bits_ftqOffset;
  wire [5:0] io_perf_0_value;
  wire [5:0] io_perf_1_value;
  wire [5:0] io_perf_2_value;
  wire [5:0] io_perf_3_value;


 DecodeStage DecodeStage(
    .clock(clock),
    .reset(reset),
    .io_redirect(io_redirect),
    .io_in_0_ready(io_in_0_ready),
    .io_in_0_valid(io_in_0_valid),
    .io_in_0_bits_instr(io_in_0_bits_instr),
    .io_in_0_bits_exceptionVec_0(io_in_0_bits_exceptionVec_0),
    .io_in_0_bits_exceptionVec_1(io_in_0_bits_exceptionVec_1),
    .io_in_0_bits_exceptionVec_2(io_in_0_bits_exceptionVec_2),
    .io_in_0_bits_exceptionVec_4(io_in_0_bits_exceptionVec_4),
    .io_in_0_bits_exceptionVec_5(io_in_0_bits_exceptionVec_5),
    .io_in_0_bits_exceptionVec_6(io_in_0_bits_exceptionVec_6),
    .io_in_0_bits_exceptionVec_7(io_in_0_bits_exceptionVec_7),
    .io_in_0_bits_exceptionVec_8(io_in_0_bits_exceptionVec_8),
    .io_in_0_bits_exceptionVec_9(io_in_0_bits_exceptionVec_9),
    .io_in_0_bits_exceptionVec_10(io_in_0_bits_exceptionVec_10),
    .io_in_0_bits_exceptionVec_11(io_in_0_bits_exceptionVec_11),
    .io_in_0_bits_exceptionVec_12(io_in_0_bits_exceptionVec_12),
    .io_in_0_bits_exceptionVec_13(io_in_0_bits_exceptionVec_13),
    .io_in_0_bits_exceptionVec_14(io_in_0_bits_exceptionVec_14),
    .io_in_0_bits_exceptionVec_15(io_in_0_bits_exceptionVec_15),
    .io_in_0_bits_exceptionVec_16(io_in_0_bits_exceptionVec_16),
    .io_in_0_bits_exceptionVec_17(io_in_0_bits_exceptionVec_17),
    .io_in_0_bits_exceptionVec_18(io_in_0_bits_exceptionVec_18),
    .io_in_0_bits_exceptionVec_19(io_in_0_bits_exceptionVec_19),
    .io_in_0_bits_exceptionVec_20(io_in_0_bits_exceptionVec_20),
    .io_in_0_bits_exceptionVec_21(io_in_0_bits_exceptionVec_21),
    .io_in_0_bits_exceptionVec_23(io_in_0_bits_exceptionVec_23),
    .io_in_0_bits_isFetchMalAddr(io_in_0_bits_isFetchMalAddr),
    .io_in_0_bits_trigger(io_in_0_bits_trigger),
    .io_in_0_bits_preDecodeInfo_isRVC(io_in_0_bits_preDecodeInfo_isRVC),
    .io_in_0_bits_preDecodeInfo_brType(io_in_0_bits_preDecodeInfo_brType),
    .io_in_0_bits_pred_taken(io_in_0_bits_pred_taken),
    .io_in_0_bits_crossPageIPFFix(io_in_0_bits_crossPageIPFFix),
    .io_in_0_bits_ftqPtr_flag(io_in_0_bits_ftqPtr_flag),
    .io_in_0_bits_ftqPtr_value(io_in_0_bits_ftqPtr_value),
    .io_in_0_bits_ftqOffset(io_in_0_bits_ftqOffset),
    .io_in_0_bits_isLastInFtqEntry(io_in_0_bits_isLastInFtqEntry),
    .io_in_1_ready(io_in_1_ready),
    .io_in_1_valid(io_in_1_valid),
    .io_in_1_bits_instr(io_in_1_bits_instr),
    .io_in_1_bits_exceptionVec_0(io_in_1_bits_exceptionVec_0),
    .io_in_1_bits_exceptionVec_1(io_in_1_bits_exceptionVec_1),
    .io_in_1_bits_exceptionVec_2(io_in_1_bits_exceptionVec_2),
    .io_in_1_bits_exceptionVec_4(io_in_1_bits_exceptionVec_4),
    .io_in_1_bits_exceptionVec_5(io_in_1_bits_exceptionVec_5),
    .io_in_1_bits_exceptionVec_6(io_in_1_bits_exceptionVec_6),
    .io_in_1_bits_exceptionVec_7(io_in_1_bits_exceptionVec_7),
    .io_in_1_bits_exceptionVec_8(io_in_1_bits_exceptionVec_8),
    .io_in_1_bits_exceptionVec_9(io_in_1_bits_exceptionVec_9),
    .io_in_1_bits_exceptionVec_10(io_in_1_bits_exceptionVec_10),
    .io_in_1_bits_exceptionVec_11(io_in_1_bits_exceptionVec_11),
    .io_in_1_bits_exceptionVec_12(io_in_1_bits_exceptionVec_12),
    .io_in_1_bits_exceptionVec_13(io_in_1_bits_exceptionVec_13),
    .io_in_1_bits_exceptionVec_14(io_in_1_bits_exceptionVec_14),
    .io_in_1_bits_exceptionVec_15(io_in_1_bits_exceptionVec_15),
    .io_in_1_bits_exceptionVec_16(io_in_1_bits_exceptionVec_16),
    .io_in_1_bits_exceptionVec_17(io_in_1_bits_exceptionVec_17),
    .io_in_1_bits_exceptionVec_18(io_in_1_bits_exceptionVec_18),
    .io_in_1_bits_exceptionVec_19(io_in_1_bits_exceptionVec_19),
    .io_in_1_bits_exceptionVec_20(io_in_1_bits_exceptionVec_20),
    .io_in_1_bits_exceptionVec_21(io_in_1_bits_exceptionVec_21),
    .io_in_1_bits_exceptionVec_23(io_in_1_bits_exceptionVec_23),
    .io_in_1_bits_isFetchMalAddr(io_in_1_bits_isFetchMalAddr),
    .io_in_1_bits_trigger(io_in_1_bits_trigger),
    .io_in_1_bits_preDecodeInfo_isRVC(io_in_1_bits_preDecodeInfo_isRVC),
    .io_in_1_bits_preDecodeInfo_brType(io_in_1_bits_preDecodeInfo_brType),
    .io_in_1_bits_pred_taken(io_in_1_bits_pred_taken),
    .io_in_1_bits_crossPageIPFFix(io_in_1_bits_crossPageIPFFix),
    .io_in_1_bits_ftqPtr_flag(io_in_1_bits_ftqPtr_flag),
    .io_in_1_bits_ftqPtr_value(io_in_1_bits_ftqPtr_value),
    .io_in_1_bits_ftqOffset(io_in_1_bits_ftqOffset),
    .io_in_1_bits_isLastInFtqEntry(io_in_1_bits_isLastInFtqEntry),
    .io_in_2_ready(io_in_2_ready),
    .io_in_2_valid(io_in_2_valid),
    .io_in_2_bits_instr(io_in_2_bits_instr),
    .io_in_2_bits_exceptionVec_0(io_in_2_bits_exceptionVec_0),
    .io_in_2_bits_exceptionVec_1(io_in_2_bits_exceptionVec_1),
    .io_in_2_bits_exceptionVec_2(io_in_2_bits_exceptionVec_2),
    .io_in_2_bits_exceptionVec_4(io_in_2_bits_exceptionVec_4),
    .io_in_2_bits_exceptionVec_5(io_in_2_bits_exceptionVec_5),
    .io_in_2_bits_exceptionVec_6(io_in_2_bits_exceptionVec_6),
    .io_in_2_bits_exceptionVec_7(io_in_2_bits_exceptionVec_7),
    .io_in_2_bits_exceptionVec_8(io_in_2_bits_exceptionVec_8),
    .io_in_2_bits_exceptionVec_9(io_in_2_bits_exceptionVec_9),
    .io_in_2_bits_exceptionVec_10(io_in_2_bits_exceptionVec_10),
    .io_in_2_bits_exceptionVec_11(io_in_2_bits_exceptionVec_11),
    .io_in_2_bits_exceptionVec_12(io_in_2_bits_exceptionVec_12),
    .io_in_2_bits_exceptionVec_13(io_in_2_bits_exceptionVec_13),
    .io_in_2_bits_exceptionVec_14(io_in_2_bits_exceptionVec_14),
    .io_in_2_bits_exceptionVec_15(io_in_2_bits_exceptionVec_15),
    .io_in_2_bits_exceptionVec_16(io_in_2_bits_exceptionVec_16),
    .io_in_2_bits_exceptionVec_17(io_in_2_bits_exceptionVec_17),
    .io_in_2_bits_exceptionVec_18(io_in_2_bits_exceptionVec_18),
    .io_in_2_bits_exceptionVec_19(io_in_2_bits_exceptionVec_19),
    .io_in_2_bits_exceptionVec_20(io_in_2_bits_exceptionVec_20),
    .io_in_2_bits_exceptionVec_21(io_in_2_bits_exceptionVec_21),
    .io_in_2_bits_exceptionVec_23(io_in_2_bits_exceptionVec_23),
    .io_in_2_bits_isFetchMalAddr(io_in_2_bits_isFetchMalAddr),
    .io_in_2_bits_trigger(io_in_2_bits_trigger),
    .io_in_2_bits_preDecodeInfo_isRVC(io_in_2_bits_preDecodeInfo_isRVC),
    .io_in_2_bits_preDecodeInfo_brType(io_in_2_bits_preDecodeInfo_brType),
    .io_in_2_bits_pred_taken(io_in_2_bits_pred_taken),
    .io_in_2_bits_crossPageIPFFix(io_in_2_bits_crossPageIPFFix),
    .io_in_2_bits_ftqPtr_flag(io_in_2_bits_ftqPtr_flag),
    .io_in_2_bits_ftqPtr_value(io_in_2_bits_ftqPtr_value),
    .io_in_2_bits_ftqOffset(io_in_2_bits_ftqOffset),
    .io_in_2_bits_isLastInFtqEntry(io_in_2_bits_isLastInFtqEntry),
    .io_in_3_ready(io_in_3_ready),
    .io_in_3_valid(io_in_3_valid),
    .io_in_3_bits_instr(io_in_3_bits_instr),
    .io_in_3_bits_exceptionVec_0(io_in_3_bits_exceptionVec_0),
    .io_in_3_bits_exceptionVec_1(io_in_3_bits_exceptionVec_1),
    .io_in_3_bits_exceptionVec_2(io_in_3_bits_exceptionVec_2),
    .io_in_3_bits_exceptionVec_4(io_in_3_bits_exceptionVec_4),
    .io_in_3_bits_exceptionVec_5(io_in_3_bits_exceptionVec_5),
    .io_in_3_bits_exceptionVec_6(io_in_3_bits_exceptionVec_6),
    .io_in_3_bits_exceptionVec_7(io_in_3_bits_exceptionVec_7),
    .io_in_3_bits_exceptionVec_8(io_in_3_bits_exceptionVec_8),
    .io_in_3_bits_exceptionVec_9(io_in_3_bits_exceptionVec_9),
    .io_in_3_bits_exceptionVec_10(io_in_3_bits_exceptionVec_10),
    .io_in_3_bits_exceptionVec_11(io_in_3_bits_exceptionVec_11),
    .io_in_3_bits_exceptionVec_12(io_in_3_bits_exceptionVec_12),
    .io_in_3_bits_exceptionVec_13(io_in_3_bits_exceptionVec_13),
    .io_in_3_bits_exceptionVec_14(io_in_3_bits_exceptionVec_14),
    .io_in_3_bits_exceptionVec_15(io_in_3_bits_exceptionVec_15),
    .io_in_3_bits_exceptionVec_16(io_in_3_bits_exceptionVec_16),
    .io_in_3_bits_exceptionVec_17(io_in_3_bits_exceptionVec_17),
    .io_in_3_bits_exceptionVec_18(io_in_3_bits_exceptionVec_18),
    .io_in_3_bits_exceptionVec_19(io_in_3_bits_exceptionVec_19),
    .io_in_3_bits_exceptionVec_20(io_in_3_bits_exceptionVec_20),
    .io_in_3_bits_exceptionVec_21(io_in_3_bits_exceptionVec_21),
    .io_in_3_bits_exceptionVec_23(io_in_3_bits_exceptionVec_23),
    .io_in_3_bits_isFetchMalAddr(io_in_3_bits_isFetchMalAddr),
    .io_in_3_bits_trigger(io_in_3_bits_trigger),
    .io_in_3_bits_preDecodeInfo_isRVC(io_in_3_bits_preDecodeInfo_isRVC),
    .io_in_3_bits_preDecodeInfo_brType(io_in_3_bits_preDecodeInfo_brType),
    .io_in_3_bits_pred_taken(io_in_3_bits_pred_taken),
    .io_in_3_bits_crossPageIPFFix(io_in_3_bits_crossPageIPFFix),
    .io_in_3_bits_ftqPtr_flag(io_in_3_bits_ftqPtr_flag),
    .io_in_3_bits_ftqPtr_value(io_in_3_bits_ftqPtr_value),
    .io_in_3_bits_ftqOffset(io_in_3_bits_ftqOffset),
    .io_in_3_bits_isLastInFtqEntry(io_in_3_bits_isLastInFtqEntry),
    .io_in_4_ready(io_in_4_ready),
    .io_in_4_valid(io_in_4_valid),
    .io_in_4_bits_instr(io_in_4_bits_instr),
    .io_in_4_bits_exceptionVec_0(io_in_4_bits_exceptionVec_0),
    .io_in_4_bits_exceptionVec_1(io_in_4_bits_exceptionVec_1),
    .io_in_4_bits_exceptionVec_2(io_in_4_bits_exceptionVec_2),
    .io_in_4_bits_exceptionVec_4(io_in_4_bits_exceptionVec_4),
    .io_in_4_bits_exceptionVec_5(io_in_4_bits_exceptionVec_5),
    .io_in_4_bits_exceptionVec_6(io_in_4_bits_exceptionVec_6),
    .io_in_4_bits_exceptionVec_7(io_in_4_bits_exceptionVec_7),
    .io_in_4_bits_exceptionVec_8(io_in_4_bits_exceptionVec_8),
    .io_in_4_bits_exceptionVec_9(io_in_4_bits_exceptionVec_9),
    .io_in_4_bits_exceptionVec_10(io_in_4_bits_exceptionVec_10),
    .io_in_4_bits_exceptionVec_11(io_in_4_bits_exceptionVec_11),
    .io_in_4_bits_exceptionVec_12(io_in_4_bits_exceptionVec_12),
    .io_in_4_bits_exceptionVec_13(io_in_4_bits_exceptionVec_13),
    .io_in_4_bits_exceptionVec_14(io_in_4_bits_exceptionVec_14),
    .io_in_4_bits_exceptionVec_15(io_in_4_bits_exceptionVec_15),
    .io_in_4_bits_exceptionVec_16(io_in_4_bits_exceptionVec_16),
    .io_in_4_bits_exceptionVec_17(io_in_4_bits_exceptionVec_17),
    .io_in_4_bits_exceptionVec_18(io_in_4_bits_exceptionVec_18),
    .io_in_4_bits_exceptionVec_19(io_in_4_bits_exceptionVec_19),
    .io_in_4_bits_exceptionVec_20(io_in_4_bits_exceptionVec_20),
    .io_in_4_bits_exceptionVec_21(io_in_4_bits_exceptionVec_21),
    .io_in_4_bits_exceptionVec_23(io_in_4_bits_exceptionVec_23),
    .io_in_4_bits_isFetchMalAddr(io_in_4_bits_isFetchMalAddr),
    .io_in_4_bits_trigger(io_in_4_bits_trigger),
    .io_in_4_bits_preDecodeInfo_isRVC(io_in_4_bits_preDecodeInfo_isRVC),
    .io_in_4_bits_preDecodeInfo_brType(io_in_4_bits_preDecodeInfo_brType),
    .io_in_4_bits_pred_taken(io_in_4_bits_pred_taken),
    .io_in_4_bits_crossPageIPFFix(io_in_4_bits_crossPageIPFFix),
    .io_in_4_bits_ftqPtr_flag(io_in_4_bits_ftqPtr_flag),
    .io_in_4_bits_ftqPtr_value(io_in_4_bits_ftqPtr_value),
    .io_in_4_bits_ftqOffset(io_in_4_bits_ftqOffset),
    .io_in_4_bits_isLastInFtqEntry(io_in_4_bits_isLastInFtqEntry),
    .io_in_5_ready(io_in_5_ready),
    .io_in_5_valid(io_in_5_valid),
    .io_in_5_bits_instr(io_in_5_bits_instr),
    .io_in_5_bits_exceptionVec_0(io_in_5_bits_exceptionVec_0),
    .io_in_5_bits_exceptionVec_1(io_in_5_bits_exceptionVec_1),
    .io_in_5_bits_exceptionVec_2(io_in_5_bits_exceptionVec_2),
    .io_in_5_bits_exceptionVec_4(io_in_5_bits_exceptionVec_4),
    .io_in_5_bits_exceptionVec_5(io_in_5_bits_exceptionVec_5),
    .io_in_5_bits_exceptionVec_6(io_in_5_bits_exceptionVec_6),
    .io_in_5_bits_exceptionVec_7(io_in_5_bits_exceptionVec_7),
    .io_in_5_bits_exceptionVec_8(io_in_5_bits_exceptionVec_8),
    .io_in_5_bits_exceptionVec_9(io_in_5_bits_exceptionVec_9),
    .io_in_5_bits_exceptionVec_10(io_in_5_bits_exceptionVec_10),
    .io_in_5_bits_exceptionVec_11(io_in_5_bits_exceptionVec_11),
    .io_in_5_bits_exceptionVec_12(io_in_5_bits_exceptionVec_12),
    .io_in_5_bits_exceptionVec_13(io_in_5_bits_exceptionVec_13),
    .io_in_5_bits_exceptionVec_14(io_in_5_bits_exceptionVec_14),
    .io_in_5_bits_exceptionVec_15(io_in_5_bits_exceptionVec_15),
    .io_in_5_bits_exceptionVec_16(io_in_5_bits_exceptionVec_16),
    .io_in_5_bits_exceptionVec_17(io_in_5_bits_exceptionVec_17),
    .io_in_5_bits_exceptionVec_18(io_in_5_bits_exceptionVec_18),
    .io_in_5_bits_exceptionVec_19(io_in_5_bits_exceptionVec_19),
    .io_in_5_bits_exceptionVec_20(io_in_5_bits_exceptionVec_20),
    .io_in_5_bits_exceptionVec_21(io_in_5_bits_exceptionVec_21),
    .io_in_5_bits_exceptionVec_23(io_in_5_bits_exceptionVec_23),
    .io_in_5_bits_isFetchMalAddr(io_in_5_bits_isFetchMalAddr),
    .io_in_5_bits_trigger(io_in_5_bits_trigger),
    .io_in_5_bits_preDecodeInfo_isRVC(io_in_5_bits_preDecodeInfo_isRVC),
    .io_in_5_bits_preDecodeInfo_brType(io_in_5_bits_preDecodeInfo_brType),
    .io_in_5_bits_pred_taken(io_in_5_bits_pred_taken),
    .io_in_5_bits_crossPageIPFFix(io_in_5_bits_crossPageIPFFix),
    .io_in_5_bits_ftqPtr_flag(io_in_5_bits_ftqPtr_flag),
    .io_in_5_bits_ftqPtr_value(io_in_5_bits_ftqPtr_value),
    .io_in_5_bits_ftqOffset(io_in_5_bits_ftqOffset),
    .io_in_5_bits_isLastInFtqEntry(io_in_5_bits_isLastInFtqEntry),
    .io_out_0_ready(io_out_0_ready),
    .io_out_0_valid(io_out_0_valid),
    .io_out_0_bits_instr(io_out_0_bits_instr),
    .io_out_0_bits_exceptionVec_0(io_out_0_bits_exceptionVec_0),
    .io_out_0_bits_exceptionVec_1(io_out_0_bits_exceptionVec_1),
    .io_out_0_bits_exceptionVec_2(io_out_0_bits_exceptionVec_2),
    .io_out_0_bits_exceptionVec_3(io_out_0_bits_exceptionVec_3),
    .io_out_0_bits_exceptionVec_4(io_out_0_bits_exceptionVec_4),
    .io_out_0_bits_exceptionVec_5(io_out_0_bits_exceptionVec_5),
    .io_out_0_bits_exceptionVec_6(io_out_0_bits_exceptionVec_6),
    .io_out_0_bits_exceptionVec_7(io_out_0_bits_exceptionVec_7),
    .io_out_0_bits_exceptionVec_8(io_out_0_bits_exceptionVec_8),
    .io_out_0_bits_exceptionVec_9(io_out_0_bits_exceptionVec_9),
    .io_out_0_bits_exceptionVec_10(io_out_0_bits_exceptionVec_10),
    .io_out_0_bits_exceptionVec_11(io_out_0_bits_exceptionVec_11),
    .io_out_0_bits_exceptionVec_12(io_out_0_bits_exceptionVec_12),
    .io_out_0_bits_exceptionVec_13(io_out_0_bits_exceptionVec_13),
    .io_out_0_bits_exceptionVec_14(io_out_0_bits_exceptionVec_14),
    .io_out_0_bits_exceptionVec_15(io_out_0_bits_exceptionVec_15),
    .io_out_0_bits_exceptionVec_16(io_out_0_bits_exceptionVec_16),
    .io_out_0_bits_exceptionVec_17(io_out_0_bits_exceptionVec_17),
    .io_out_0_bits_exceptionVec_18(io_out_0_bits_exceptionVec_18),
    .io_out_0_bits_exceptionVec_19(io_out_0_bits_exceptionVec_19),
    .io_out_0_bits_exceptionVec_20(io_out_0_bits_exceptionVec_20),
    .io_out_0_bits_exceptionVec_21(io_out_0_bits_exceptionVec_21),
    .io_out_0_bits_exceptionVec_22(io_out_0_bits_exceptionVec_22),
    .io_out_0_bits_exceptionVec_23(io_out_0_bits_exceptionVec_23),
    .io_out_0_bits_isFetchMalAddr(io_out_0_bits_isFetchMalAddr),
    .io_out_0_bits_trigger(io_out_0_bits_trigger),
    .io_out_0_bits_preDecodeInfo_isRVC(io_out_0_bits_preDecodeInfo_isRVC),
    .io_out_0_bits_preDecodeInfo_brType(io_out_0_bits_preDecodeInfo_brType),
    .io_out_0_bits_pred_taken(io_out_0_bits_pred_taken),
    .io_out_0_bits_crossPageIPFFix(io_out_0_bits_crossPageIPFFix),
    .io_out_0_bits_ftqPtr_flag(io_out_0_bits_ftqPtr_flag),
    .io_out_0_bits_ftqPtr_value(io_out_0_bits_ftqPtr_value),
    .io_out_0_bits_ftqOffset(io_out_0_bits_ftqOffset),
    .io_out_0_bits_srcType_0(io_out_0_bits_srcType_0),
    .io_out_0_bits_srcType_1(io_out_0_bits_srcType_1),
    .io_out_0_bits_srcType_2(io_out_0_bits_srcType_2),
    .io_out_0_bits_srcType_3(io_out_0_bits_srcType_3),
    .io_out_0_bits_srcType_4(io_out_0_bits_srcType_4),
    .io_out_0_bits_lsrc_0(io_out_0_bits_lsrc_0),
    .io_out_0_bits_lsrc_1(io_out_0_bits_lsrc_1),
    .io_out_0_bits_lsrc_2(io_out_0_bits_lsrc_2),
    .io_out_0_bits_ldest(io_out_0_bits_ldest),
    .io_out_0_bits_fuType(io_out_0_bits_fuType),
    .io_out_0_bits_fuOpType(io_out_0_bits_fuOpType),
    .io_out_0_bits_rfWen(io_out_0_bits_rfWen),
    .io_out_0_bits_fpWen(io_out_0_bits_fpWen),
    .io_out_0_bits_vecWen(io_out_0_bits_vecWen),
    .io_out_0_bits_v0Wen(io_out_0_bits_v0Wen),
    .io_out_0_bits_vlWen(io_out_0_bits_vlWen),
    .io_out_0_bits_isXSTrap(io_out_0_bits_isXSTrap),
    .io_out_0_bits_waitForward(io_out_0_bits_waitForward),
    .io_out_0_bits_blockBackward(io_out_0_bits_blockBackward),
    .io_out_0_bits_flushPipe(io_out_0_bits_flushPipe),
    .io_out_0_bits_canRobCompress(io_out_0_bits_canRobCompress),
    .io_out_0_bits_selImm(io_out_0_bits_selImm),
    .io_out_0_bits_imm(io_out_0_bits_imm),
    .io_out_0_bits_fpu_typeTagOut(io_out_0_bits_fpu_typeTagOut),
    .io_out_0_bits_fpu_wflags(io_out_0_bits_fpu_wflags),
    .io_out_0_bits_fpu_typ(io_out_0_bits_fpu_typ),
    .io_out_0_bits_fpu_fmt(io_out_0_bits_fpu_fmt),
    .io_out_0_bits_fpu_rm(io_out_0_bits_fpu_rm),
    .io_out_0_bits_vpu_vill(io_out_0_bits_vpu_vill),
    .io_out_0_bits_vpu_vma(io_out_0_bits_vpu_vma),
    .io_out_0_bits_vpu_vta(io_out_0_bits_vpu_vta),
    .io_out_0_bits_vpu_vsew(io_out_0_bits_vpu_vsew),
    .io_out_0_bits_vpu_vlmul(io_out_0_bits_vpu_vlmul),
    .io_out_0_bits_vpu_specVill(io_out_0_bits_vpu_specVill),
    .io_out_0_bits_vpu_specVma(io_out_0_bits_vpu_specVma),
    .io_out_0_bits_vpu_specVta(io_out_0_bits_vpu_specVta),
    .io_out_0_bits_vpu_specVsew(io_out_0_bits_vpu_specVsew),
    .io_out_0_bits_vpu_specVlmul(io_out_0_bits_vpu_specVlmul),
    .io_out_0_bits_vpu_vm(io_out_0_bits_vpu_vm),
    .io_out_0_bits_vpu_vstart(io_out_0_bits_vpu_vstart),
    .io_out_0_bits_vpu_fpu_isFoldTo1_2(io_out_0_bits_vpu_fpu_isFoldTo1_2),
    .io_out_0_bits_vpu_fpu_isFoldTo1_4(io_out_0_bits_vpu_fpu_isFoldTo1_4),
    .io_out_0_bits_vpu_fpu_isFoldTo1_8(io_out_0_bits_vpu_fpu_isFoldTo1_8),
    .io_out_0_bits_vpu_nf(io_out_0_bits_vpu_nf),
    .io_out_0_bits_vpu_veew(io_out_0_bits_vpu_veew),
    .io_out_0_bits_vpu_isExt(io_out_0_bits_vpu_isExt),
    .io_out_0_bits_vpu_isNarrow(io_out_0_bits_vpu_isNarrow),
    .io_out_0_bits_vpu_isDstMask(io_out_0_bits_vpu_isDstMask),
    .io_out_0_bits_vpu_isOpMask(io_out_0_bits_vpu_isOpMask),
    .io_out_0_bits_vpu_isDependOldVd(io_out_0_bits_vpu_isDependOldVd),
    .io_out_0_bits_vpu_isWritePartVd(io_out_0_bits_vpu_isWritePartVd),
    .io_out_0_bits_vpu_isVleff(io_out_0_bits_vpu_isVleff),
    .io_out_0_bits_vlsInstr(io_out_0_bits_vlsInstr),
    .io_out_0_bits_wfflags(io_out_0_bits_wfflags),
    .io_out_0_bits_isMove(io_out_0_bits_isMove),
    .io_out_0_bits_uopIdx(io_out_0_bits_uopIdx),
    .io_out_0_bits_uopSplitType(io_out_0_bits_uopSplitType),
    .io_out_0_bits_isVset(io_out_0_bits_isVset),
    .io_out_0_bits_firstUop(io_out_0_bits_firstUop),
    .io_out_0_bits_lastUop(io_out_0_bits_lastUop),
    .io_out_0_bits_numWB(io_out_0_bits_numWB),
    .io_out_0_bits_commitType(io_out_0_bits_commitType),
    .io_out_1_ready(io_out_1_ready),
    .io_out_1_valid(io_out_1_valid),
    .io_out_1_bits_instr(io_out_1_bits_instr),
    .io_out_1_bits_exceptionVec_0(io_out_1_bits_exceptionVec_0),
    .io_out_1_bits_exceptionVec_1(io_out_1_bits_exceptionVec_1),
    .io_out_1_bits_exceptionVec_2(io_out_1_bits_exceptionVec_2),
    .io_out_1_bits_exceptionVec_3(io_out_1_bits_exceptionVec_3),
    .io_out_1_bits_exceptionVec_4(io_out_1_bits_exceptionVec_4),
    .io_out_1_bits_exceptionVec_5(io_out_1_bits_exceptionVec_5),
    .io_out_1_bits_exceptionVec_6(io_out_1_bits_exceptionVec_6),
    .io_out_1_bits_exceptionVec_7(io_out_1_bits_exceptionVec_7),
    .io_out_1_bits_exceptionVec_8(io_out_1_bits_exceptionVec_8),
    .io_out_1_bits_exceptionVec_9(io_out_1_bits_exceptionVec_9),
    .io_out_1_bits_exceptionVec_10(io_out_1_bits_exceptionVec_10),
    .io_out_1_bits_exceptionVec_11(io_out_1_bits_exceptionVec_11),
    .io_out_1_bits_exceptionVec_12(io_out_1_bits_exceptionVec_12),
    .io_out_1_bits_exceptionVec_13(io_out_1_bits_exceptionVec_13),
    .io_out_1_bits_exceptionVec_14(io_out_1_bits_exceptionVec_14),
    .io_out_1_bits_exceptionVec_15(io_out_1_bits_exceptionVec_15),
    .io_out_1_bits_exceptionVec_16(io_out_1_bits_exceptionVec_16),
    .io_out_1_bits_exceptionVec_17(io_out_1_bits_exceptionVec_17),
    .io_out_1_bits_exceptionVec_18(io_out_1_bits_exceptionVec_18),
    .io_out_1_bits_exceptionVec_19(io_out_1_bits_exceptionVec_19),
    .io_out_1_bits_exceptionVec_20(io_out_1_bits_exceptionVec_20),
    .io_out_1_bits_exceptionVec_21(io_out_1_bits_exceptionVec_21),
    .io_out_1_bits_exceptionVec_22(io_out_1_bits_exceptionVec_22),
    .io_out_1_bits_exceptionVec_23(io_out_1_bits_exceptionVec_23),
    .io_out_1_bits_isFetchMalAddr(io_out_1_bits_isFetchMalAddr),
    .io_out_1_bits_trigger(io_out_1_bits_trigger),
    .io_out_1_bits_preDecodeInfo_isRVC(io_out_1_bits_preDecodeInfo_isRVC),
    .io_out_1_bits_preDecodeInfo_brType(io_out_1_bits_preDecodeInfo_brType),
    .io_out_1_bits_pred_taken(io_out_1_bits_pred_taken),
    .io_out_1_bits_crossPageIPFFix(io_out_1_bits_crossPageIPFFix),
    .io_out_1_bits_ftqPtr_flag(io_out_1_bits_ftqPtr_flag),
    .io_out_1_bits_ftqPtr_value(io_out_1_bits_ftqPtr_value),
    .io_out_1_bits_ftqOffset(io_out_1_bits_ftqOffset),
    .io_out_1_bits_srcType_0(io_out_1_bits_srcType_0),
    .io_out_1_bits_srcType_1(io_out_1_bits_srcType_1),
    .io_out_1_bits_srcType_2(io_out_1_bits_srcType_2),
    .io_out_1_bits_srcType_3(io_out_1_bits_srcType_3),
    .io_out_1_bits_srcType_4(io_out_1_bits_srcType_4),
    .io_out_1_bits_lsrc_0(io_out_1_bits_lsrc_0),
    .io_out_1_bits_lsrc_1(io_out_1_bits_lsrc_1),
    .io_out_1_bits_lsrc_2(io_out_1_bits_lsrc_2),
    .io_out_1_bits_ldest(io_out_1_bits_ldest),
    .io_out_1_bits_fuType(io_out_1_bits_fuType),
    .io_out_1_bits_fuOpType(io_out_1_bits_fuOpType),
    .io_out_1_bits_rfWen(io_out_1_bits_rfWen),
    .io_out_1_bits_fpWen(io_out_1_bits_fpWen),
    .io_out_1_bits_vecWen(io_out_1_bits_vecWen),
    .io_out_1_bits_v0Wen(io_out_1_bits_v0Wen),
    .io_out_1_bits_vlWen(io_out_1_bits_vlWen),
    .io_out_1_bits_isXSTrap(io_out_1_bits_isXSTrap),
    .io_out_1_bits_waitForward(io_out_1_bits_waitForward),
    .io_out_1_bits_blockBackward(io_out_1_bits_blockBackward),
    .io_out_1_bits_flushPipe(io_out_1_bits_flushPipe),
    .io_out_1_bits_canRobCompress(io_out_1_bits_canRobCompress),
    .io_out_1_bits_selImm(io_out_1_bits_selImm),
    .io_out_1_bits_imm(io_out_1_bits_imm),
    .io_out_1_bits_fpu_typeTagOut(io_out_1_bits_fpu_typeTagOut),
    .io_out_1_bits_fpu_wflags(io_out_1_bits_fpu_wflags),
    .io_out_1_bits_fpu_typ(io_out_1_bits_fpu_typ),
    .io_out_1_bits_fpu_fmt(io_out_1_bits_fpu_fmt),
    .io_out_1_bits_fpu_rm(io_out_1_bits_fpu_rm),
    .io_out_1_bits_vpu_vill(io_out_1_bits_vpu_vill),
    .io_out_1_bits_vpu_vma(io_out_1_bits_vpu_vma),
    .io_out_1_bits_vpu_vta(io_out_1_bits_vpu_vta),
    .io_out_1_bits_vpu_vsew(io_out_1_bits_vpu_vsew),
    .io_out_1_bits_vpu_vlmul(io_out_1_bits_vpu_vlmul),
    .io_out_1_bits_vpu_specVill(io_out_1_bits_vpu_specVill),
    .io_out_1_bits_vpu_specVma(io_out_1_bits_vpu_specVma),
    .io_out_1_bits_vpu_specVta(io_out_1_bits_vpu_specVta),
    .io_out_1_bits_vpu_specVsew(io_out_1_bits_vpu_specVsew),
    .io_out_1_bits_vpu_specVlmul(io_out_1_bits_vpu_specVlmul),
    .io_out_1_bits_vpu_vm(io_out_1_bits_vpu_vm),
    .io_out_1_bits_vpu_vstart(io_out_1_bits_vpu_vstart),
    .io_out_1_bits_vpu_fpu_isFoldTo1_2(io_out_1_bits_vpu_fpu_isFoldTo1_2),
    .io_out_1_bits_vpu_fpu_isFoldTo1_4(io_out_1_bits_vpu_fpu_isFoldTo1_4),
    .io_out_1_bits_vpu_fpu_isFoldTo1_8(io_out_1_bits_vpu_fpu_isFoldTo1_8),
    .io_out_1_bits_vpu_nf(io_out_1_bits_vpu_nf),
    .io_out_1_bits_vpu_veew(io_out_1_bits_vpu_veew),
    .io_out_1_bits_vpu_isExt(io_out_1_bits_vpu_isExt),
    .io_out_1_bits_vpu_isNarrow(io_out_1_bits_vpu_isNarrow),
    .io_out_1_bits_vpu_isDstMask(io_out_1_bits_vpu_isDstMask),
    .io_out_1_bits_vpu_isOpMask(io_out_1_bits_vpu_isOpMask),
    .io_out_1_bits_vpu_isDependOldVd(io_out_1_bits_vpu_isDependOldVd),
    .io_out_1_bits_vpu_isWritePartVd(io_out_1_bits_vpu_isWritePartVd),
    .io_out_1_bits_vpu_isVleff(io_out_1_bits_vpu_isVleff),
    .io_out_1_bits_vlsInstr(io_out_1_bits_vlsInstr),
    .io_out_1_bits_wfflags(io_out_1_bits_wfflags),
    .io_out_1_bits_isMove(io_out_1_bits_isMove),
    .io_out_1_bits_uopIdx(io_out_1_bits_uopIdx),
    .io_out_1_bits_uopSplitType(io_out_1_bits_uopSplitType),
    .io_out_1_bits_isVset(io_out_1_bits_isVset),
    .io_out_1_bits_firstUop(io_out_1_bits_firstUop),
    .io_out_1_bits_lastUop(io_out_1_bits_lastUop),
    .io_out_1_bits_numWB(io_out_1_bits_numWB),
    .io_out_1_bits_commitType(io_out_1_bits_commitType),
    .io_out_2_ready(io_out_2_ready),
    .io_out_2_valid(io_out_2_valid),
    .io_out_2_bits_instr(io_out_2_bits_instr),
    .io_out_2_bits_exceptionVec_0(io_out_2_bits_exceptionVec_0),
    .io_out_2_bits_exceptionVec_1(io_out_2_bits_exceptionVec_1),
    .io_out_2_bits_exceptionVec_2(io_out_2_bits_exceptionVec_2),
    .io_out_2_bits_exceptionVec_3(io_out_2_bits_exceptionVec_3),
    .io_out_2_bits_exceptionVec_4(io_out_2_bits_exceptionVec_4),
    .io_out_2_bits_exceptionVec_5(io_out_2_bits_exceptionVec_5),
    .io_out_2_bits_exceptionVec_6(io_out_2_bits_exceptionVec_6),
    .io_out_2_bits_exceptionVec_7(io_out_2_bits_exceptionVec_7),
    .io_out_2_bits_exceptionVec_8(io_out_2_bits_exceptionVec_8),
    .io_out_2_bits_exceptionVec_9(io_out_2_bits_exceptionVec_9),
    .io_out_2_bits_exceptionVec_10(io_out_2_bits_exceptionVec_10),
    .io_out_2_bits_exceptionVec_11(io_out_2_bits_exceptionVec_11),
    .io_out_2_bits_exceptionVec_12(io_out_2_bits_exceptionVec_12),
    .io_out_2_bits_exceptionVec_13(io_out_2_bits_exceptionVec_13),
    .io_out_2_bits_exceptionVec_14(io_out_2_bits_exceptionVec_14),
    .io_out_2_bits_exceptionVec_15(io_out_2_bits_exceptionVec_15),
    .io_out_2_bits_exceptionVec_16(io_out_2_bits_exceptionVec_16),
    .io_out_2_bits_exceptionVec_17(io_out_2_bits_exceptionVec_17),
    .io_out_2_bits_exceptionVec_18(io_out_2_bits_exceptionVec_18),
    .io_out_2_bits_exceptionVec_19(io_out_2_bits_exceptionVec_19),
    .io_out_2_bits_exceptionVec_20(io_out_2_bits_exceptionVec_20),
    .io_out_2_bits_exceptionVec_21(io_out_2_bits_exceptionVec_21),
    .io_out_2_bits_exceptionVec_22(io_out_2_bits_exceptionVec_22),
    .io_out_2_bits_exceptionVec_23(io_out_2_bits_exceptionVec_23),
    .io_out_2_bits_isFetchMalAddr(io_out_2_bits_isFetchMalAddr),
    .io_out_2_bits_trigger(io_out_2_bits_trigger),
    .io_out_2_bits_preDecodeInfo_isRVC(io_out_2_bits_preDecodeInfo_isRVC),
    .io_out_2_bits_preDecodeInfo_brType(io_out_2_bits_preDecodeInfo_brType),
    .io_out_2_bits_pred_taken(io_out_2_bits_pred_taken),
    .io_out_2_bits_crossPageIPFFix(io_out_2_bits_crossPageIPFFix),
    .io_out_2_bits_ftqPtr_flag(io_out_2_bits_ftqPtr_flag),
    .io_out_2_bits_ftqPtr_value(io_out_2_bits_ftqPtr_value),
    .io_out_2_bits_ftqOffset(io_out_2_bits_ftqOffset),
    .io_out_2_bits_srcType_0(io_out_2_bits_srcType_0),
    .io_out_2_bits_srcType_1(io_out_2_bits_srcType_1),
    .io_out_2_bits_srcType_2(io_out_2_bits_srcType_2),
    .io_out_2_bits_srcType_3(io_out_2_bits_srcType_3),
    .io_out_2_bits_srcType_4(io_out_2_bits_srcType_4),
    .io_out_2_bits_lsrc_0(io_out_2_bits_lsrc_0),
    .io_out_2_bits_lsrc_1(io_out_2_bits_lsrc_1),
    .io_out_2_bits_lsrc_2(io_out_2_bits_lsrc_2),
    .io_out_2_bits_ldest(io_out_2_bits_ldest),
    .io_out_2_bits_fuType(io_out_2_bits_fuType),
    .io_out_2_bits_fuOpType(io_out_2_bits_fuOpType),
    .io_out_2_bits_rfWen(io_out_2_bits_rfWen),
    .io_out_2_bits_fpWen(io_out_2_bits_fpWen),
    .io_out_2_bits_vecWen(io_out_2_bits_vecWen),
    .io_out_2_bits_v0Wen(io_out_2_bits_v0Wen),
    .io_out_2_bits_vlWen(io_out_2_bits_vlWen),
    .io_out_2_bits_isXSTrap(io_out_2_bits_isXSTrap),
    .io_out_2_bits_waitForward(io_out_2_bits_waitForward),
    .io_out_2_bits_blockBackward(io_out_2_bits_blockBackward),
    .io_out_2_bits_flushPipe(io_out_2_bits_flushPipe),
    .io_out_2_bits_canRobCompress(io_out_2_bits_canRobCompress),
    .io_out_2_bits_selImm(io_out_2_bits_selImm),
    .io_out_2_bits_imm(io_out_2_bits_imm),
    .io_out_2_bits_fpu_typeTagOut(io_out_2_bits_fpu_typeTagOut),
    .io_out_2_bits_fpu_wflags(io_out_2_bits_fpu_wflags),
    .io_out_2_bits_fpu_typ(io_out_2_bits_fpu_typ),
    .io_out_2_bits_fpu_fmt(io_out_2_bits_fpu_fmt),
    .io_out_2_bits_fpu_rm(io_out_2_bits_fpu_rm),
    .io_out_2_bits_vpu_vill(io_out_2_bits_vpu_vill),
    .io_out_2_bits_vpu_vma(io_out_2_bits_vpu_vma),
    .io_out_2_bits_vpu_vta(io_out_2_bits_vpu_vta),
    .io_out_2_bits_vpu_vsew(io_out_2_bits_vpu_vsew),
    .io_out_2_bits_vpu_vlmul(io_out_2_bits_vpu_vlmul),
    .io_out_2_bits_vpu_specVill(io_out_2_bits_vpu_specVill),
    .io_out_2_bits_vpu_specVma(io_out_2_bits_vpu_specVma),
    .io_out_2_bits_vpu_specVta(io_out_2_bits_vpu_specVta),
    .io_out_2_bits_vpu_specVsew(io_out_2_bits_vpu_specVsew),
    .io_out_2_bits_vpu_specVlmul(io_out_2_bits_vpu_specVlmul),
    .io_out_2_bits_vpu_vm(io_out_2_bits_vpu_vm),
    .io_out_2_bits_vpu_vstart(io_out_2_bits_vpu_vstart),
    .io_out_2_bits_vpu_fpu_isFoldTo1_2(io_out_2_bits_vpu_fpu_isFoldTo1_2),
    .io_out_2_bits_vpu_fpu_isFoldTo1_4(io_out_2_bits_vpu_fpu_isFoldTo1_4),
    .io_out_2_bits_vpu_fpu_isFoldTo1_8(io_out_2_bits_vpu_fpu_isFoldTo1_8),
    .io_out_2_bits_vpu_nf(io_out_2_bits_vpu_nf),
    .io_out_2_bits_vpu_veew(io_out_2_bits_vpu_veew),
    .io_out_2_bits_vpu_isExt(io_out_2_bits_vpu_isExt),
    .io_out_2_bits_vpu_isNarrow(io_out_2_bits_vpu_isNarrow),
    .io_out_2_bits_vpu_isDstMask(io_out_2_bits_vpu_isDstMask),
    .io_out_2_bits_vpu_isOpMask(io_out_2_bits_vpu_isOpMask),
    .io_out_2_bits_vpu_isDependOldVd(io_out_2_bits_vpu_isDependOldVd),
    .io_out_2_bits_vpu_isWritePartVd(io_out_2_bits_vpu_isWritePartVd),
    .io_out_2_bits_vpu_isVleff(io_out_2_bits_vpu_isVleff),
    .io_out_2_bits_vlsInstr(io_out_2_bits_vlsInstr),
    .io_out_2_bits_wfflags(io_out_2_bits_wfflags),
    .io_out_2_bits_isMove(io_out_2_bits_isMove),
    .io_out_2_bits_uopIdx(io_out_2_bits_uopIdx),
    .io_out_2_bits_uopSplitType(io_out_2_bits_uopSplitType),
    .io_out_2_bits_isVset(io_out_2_bits_isVset),
    .io_out_2_bits_firstUop(io_out_2_bits_firstUop),
    .io_out_2_bits_lastUop(io_out_2_bits_lastUop),
    .io_out_2_bits_numWB(io_out_2_bits_numWB),
    .io_out_2_bits_commitType(io_out_2_bits_commitType),
    .io_out_3_ready(io_out_3_ready),
    .io_out_3_valid(io_out_3_valid),
    .io_out_3_bits_instr(io_out_3_bits_instr),
    .io_out_3_bits_exceptionVec_0(io_out_3_bits_exceptionVec_0),
    .io_out_3_bits_exceptionVec_1(io_out_3_bits_exceptionVec_1),
    .io_out_3_bits_exceptionVec_2(io_out_3_bits_exceptionVec_2),
    .io_out_3_bits_exceptionVec_3(io_out_3_bits_exceptionVec_3),
    .io_out_3_bits_exceptionVec_4(io_out_3_bits_exceptionVec_4),
    .io_out_3_bits_exceptionVec_5(io_out_3_bits_exceptionVec_5),
    .io_out_3_bits_exceptionVec_6(io_out_3_bits_exceptionVec_6),
    .io_out_3_bits_exceptionVec_7(io_out_3_bits_exceptionVec_7),
    .io_out_3_bits_exceptionVec_8(io_out_3_bits_exceptionVec_8),
    .io_out_3_bits_exceptionVec_9(io_out_3_bits_exceptionVec_9),
    .io_out_3_bits_exceptionVec_10(io_out_3_bits_exceptionVec_10),
    .io_out_3_bits_exceptionVec_11(io_out_3_bits_exceptionVec_11),
    .io_out_3_bits_exceptionVec_12(io_out_3_bits_exceptionVec_12),
    .io_out_3_bits_exceptionVec_13(io_out_3_bits_exceptionVec_13),
    .io_out_3_bits_exceptionVec_14(io_out_3_bits_exceptionVec_14),
    .io_out_3_bits_exceptionVec_15(io_out_3_bits_exceptionVec_15),
    .io_out_3_bits_exceptionVec_16(io_out_3_bits_exceptionVec_16),
    .io_out_3_bits_exceptionVec_17(io_out_3_bits_exceptionVec_17),
    .io_out_3_bits_exceptionVec_18(io_out_3_bits_exceptionVec_18),
    .io_out_3_bits_exceptionVec_19(io_out_3_bits_exceptionVec_19),
    .io_out_3_bits_exceptionVec_20(io_out_3_bits_exceptionVec_20),
    .io_out_3_bits_exceptionVec_21(io_out_3_bits_exceptionVec_21),
    .io_out_3_bits_exceptionVec_22(io_out_3_bits_exceptionVec_22),
    .io_out_3_bits_exceptionVec_23(io_out_3_bits_exceptionVec_23),
    .io_out_3_bits_isFetchMalAddr(io_out_3_bits_isFetchMalAddr),
    .io_out_3_bits_trigger(io_out_3_bits_trigger),
    .io_out_3_bits_preDecodeInfo_isRVC(io_out_3_bits_preDecodeInfo_isRVC),
    .io_out_3_bits_preDecodeInfo_brType(io_out_3_bits_preDecodeInfo_brType),
    .io_out_3_bits_pred_taken(io_out_3_bits_pred_taken),
    .io_out_3_bits_crossPageIPFFix(io_out_3_bits_crossPageIPFFix),
    .io_out_3_bits_ftqPtr_flag(io_out_3_bits_ftqPtr_flag),
    .io_out_3_bits_ftqPtr_value(io_out_3_bits_ftqPtr_value),
    .io_out_3_bits_ftqOffset(io_out_3_bits_ftqOffset),
    .io_out_3_bits_srcType_0(io_out_3_bits_srcType_0),
    .io_out_3_bits_srcType_1(io_out_3_bits_srcType_1),
    .io_out_3_bits_srcType_2(io_out_3_bits_srcType_2),
    .io_out_3_bits_srcType_3(io_out_3_bits_srcType_3),
    .io_out_3_bits_srcType_4(io_out_3_bits_srcType_4),
    .io_out_3_bits_lsrc_0(io_out_3_bits_lsrc_0),
    .io_out_3_bits_lsrc_1(io_out_3_bits_lsrc_1),
    .io_out_3_bits_lsrc_2(io_out_3_bits_lsrc_2),
    .io_out_3_bits_ldest(io_out_3_bits_ldest),
    .io_out_3_bits_fuType(io_out_3_bits_fuType),
    .io_out_3_bits_fuOpType(io_out_3_bits_fuOpType),
    .io_out_3_bits_rfWen(io_out_3_bits_rfWen),
    .io_out_3_bits_fpWen(io_out_3_bits_fpWen),
    .io_out_3_bits_vecWen(io_out_3_bits_vecWen),
    .io_out_3_bits_v0Wen(io_out_3_bits_v0Wen),
    .io_out_3_bits_vlWen(io_out_3_bits_vlWen),
    .io_out_3_bits_isXSTrap(io_out_3_bits_isXSTrap),
    .io_out_3_bits_waitForward(io_out_3_bits_waitForward),
    .io_out_3_bits_blockBackward(io_out_3_bits_blockBackward),
    .io_out_3_bits_flushPipe(io_out_3_bits_flushPipe),
    .io_out_3_bits_canRobCompress(io_out_3_bits_canRobCompress),
    .io_out_3_bits_selImm(io_out_3_bits_selImm),
    .io_out_3_bits_imm(io_out_3_bits_imm),
    .io_out_3_bits_fpu_typeTagOut(io_out_3_bits_fpu_typeTagOut),
    .io_out_3_bits_fpu_wflags(io_out_3_bits_fpu_wflags),
    .io_out_3_bits_fpu_typ(io_out_3_bits_fpu_typ),
    .io_out_3_bits_fpu_fmt(io_out_3_bits_fpu_fmt),
    .io_out_3_bits_fpu_rm(io_out_3_bits_fpu_rm),
    .io_out_3_bits_vpu_vill(io_out_3_bits_vpu_vill),
    .io_out_3_bits_vpu_vma(io_out_3_bits_vpu_vma),
    .io_out_3_bits_vpu_vta(io_out_3_bits_vpu_vta),
    .io_out_3_bits_vpu_vsew(io_out_3_bits_vpu_vsew),
    .io_out_3_bits_vpu_vlmul(io_out_3_bits_vpu_vlmul),
    .io_out_3_bits_vpu_specVill(io_out_3_bits_vpu_specVill),
    .io_out_3_bits_vpu_specVma(io_out_3_bits_vpu_specVma),
    .io_out_3_bits_vpu_specVta(io_out_3_bits_vpu_specVta),
    .io_out_3_bits_vpu_specVsew(io_out_3_bits_vpu_specVsew),
    .io_out_3_bits_vpu_specVlmul(io_out_3_bits_vpu_specVlmul),
    .io_out_3_bits_vpu_vm(io_out_3_bits_vpu_vm),
    .io_out_3_bits_vpu_vstart(io_out_3_bits_vpu_vstart),
    .io_out_3_bits_vpu_fpu_isFoldTo1_2(io_out_3_bits_vpu_fpu_isFoldTo1_2),
    .io_out_3_bits_vpu_fpu_isFoldTo1_4(io_out_3_bits_vpu_fpu_isFoldTo1_4),
    .io_out_3_bits_vpu_fpu_isFoldTo1_8(io_out_3_bits_vpu_fpu_isFoldTo1_8),
    .io_out_3_bits_vpu_nf(io_out_3_bits_vpu_nf),
    .io_out_3_bits_vpu_veew(io_out_3_bits_vpu_veew),
    .io_out_3_bits_vpu_isExt(io_out_3_bits_vpu_isExt),
    .io_out_3_bits_vpu_isNarrow(io_out_3_bits_vpu_isNarrow),
    .io_out_3_bits_vpu_isDstMask(io_out_3_bits_vpu_isDstMask),
    .io_out_3_bits_vpu_isOpMask(io_out_3_bits_vpu_isOpMask),
    .io_out_3_bits_vpu_isDependOldVd(io_out_3_bits_vpu_isDependOldVd),
    .io_out_3_bits_vpu_isWritePartVd(io_out_3_bits_vpu_isWritePartVd),
    .io_out_3_bits_vpu_isVleff(io_out_3_bits_vpu_isVleff),
    .io_out_3_bits_vlsInstr(io_out_3_bits_vlsInstr),
    .io_out_3_bits_wfflags(io_out_3_bits_wfflags),
    .io_out_3_bits_isMove(io_out_3_bits_isMove),
    .io_out_3_bits_uopIdx(io_out_3_bits_uopIdx),
    .io_out_3_bits_uopSplitType(io_out_3_bits_uopSplitType),
    .io_out_3_bits_isVset(io_out_3_bits_isVset),
    .io_out_3_bits_firstUop(io_out_3_bits_firstUop),
    .io_out_3_bits_lastUop(io_out_3_bits_lastUop),
    .io_out_3_bits_numWB(io_out_3_bits_numWB),
    .io_out_3_bits_commitType(io_out_3_bits_commitType),
    .io_out_4_ready(io_out_4_ready),
    .io_out_4_valid(io_out_4_valid),
    .io_out_4_bits_instr(io_out_4_bits_instr),
    .io_out_4_bits_exceptionVec_0(io_out_4_bits_exceptionVec_0),
    .io_out_4_bits_exceptionVec_1(io_out_4_bits_exceptionVec_1),
    .io_out_4_bits_exceptionVec_2(io_out_4_bits_exceptionVec_2),
    .io_out_4_bits_exceptionVec_3(io_out_4_bits_exceptionVec_3),
    .io_out_4_bits_exceptionVec_4(io_out_4_bits_exceptionVec_4),
    .io_out_4_bits_exceptionVec_5(io_out_4_bits_exceptionVec_5),
    .io_out_4_bits_exceptionVec_6(io_out_4_bits_exceptionVec_6),
    .io_out_4_bits_exceptionVec_7(io_out_4_bits_exceptionVec_7),
    .io_out_4_bits_exceptionVec_8(io_out_4_bits_exceptionVec_8),
    .io_out_4_bits_exceptionVec_9(io_out_4_bits_exceptionVec_9),
    .io_out_4_bits_exceptionVec_10(io_out_4_bits_exceptionVec_10),
    .io_out_4_bits_exceptionVec_11(io_out_4_bits_exceptionVec_11),
    .io_out_4_bits_exceptionVec_12(io_out_4_bits_exceptionVec_12),
    .io_out_4_bits_exceptionVec_13(io_out_4_bits_exceptionVec_13),
    .io_out_4_bits_exceptionVec_14(io_out_4_bits_exceptionVec_14),
    .io_out_4_bits_exceptionVec_15(io_out_4_bits_exceptionVec_15),
    .io_out_4_bits_exceptionVec_16(io_out_4_bits_exceptionVec_16),
    .io_out_4_bits_exceptionVec_17(io_out_4_bits_exceptionVec_17),
    .io_out_4_bits_exceptionVec_18(io_out_4_bits_exceptionVec_18),
    .io_out_4_bits_exceptionVec_19(io_out_4_bits_exceptionVec_19),
    .io_out_4_bits_exceptionVec_20(io_out_4_bits_exceptionVec_20),
    .io_out_4_bits_exceptionVec_21(io_out_4_bits_exceptionVec_21),
    .io_out_4_bits_exceptionVec_22(io_out_4_bits_exceptionVec_22),
    .io_out_4_bits_exceptionVec_23(io_out_4_bits_exceptionVec_23),
    .io_out_4_bits_isFetchMalAddr(io_out_4_bits_isFetchMalAddr),
    .io_out_4_bits_trigger(io_out_4_bits_trigger),
    .io_out_4_bits_preDecodeInfo_isRVC(io_out_4_bits_preDecodeInfo_isRVC),
    .io_out_4_bits_preDecodeInfo_brType(io_out_4_bits_preDecodeInfo_brType),
    .io_out_4_bits_pred_taken(io_out_4_bits_pred_taken),
    .io_out_4_bits_crossPageIPFFix(io_out_4_bits_crossPageIPFFix),
    .io_out_4_bits_ftqPtr_flag(io_out_4_bits_ftqPtr_flag),
    .io_out_4_bits_ftqPtr_value(io_out_4_bits_ftqPtr_value),
    .io_out_4_bits_ftqOffset(io_out_4_bits_ftqOffset),
    .io_out_4_bits_srcType_0(io_out_4_bits_srcType_0),
    .io_out_4_bits_srcType_1(io_out_4_bits_srcType_1),
    .io_out_4_bits_srcType_2(io_out_4_bits_srcType_2),
    .io_out_4_bits_srcType_3(io_out_4_bits_srcType_3),
    .io_out_4_bits_srcType_4(io_out_4_bits_srcType_4),
    .io_out_4_bits_lsrc_0(io_out_4_bits_lsrc_0),
    .io_out_4_bits_lsrc_1(io_out_4_bits_lsrc_1),
    .io_out_4_bits_lsrc_2(io_out_4_bits_lsrc_2),
    .io_out_4_bits_ldest(io_out_4_bits_ldest),
    .io_out_4_bits_fuType(io_out_4_bits_fuType),
    .io_out_4_bits_fuOpType(io_out_4_bits_fuOpType),
    .io_out_4_bits_rfWen(io_out_4_bits_rfWen),
    .io_out_4_bits_fpWen(io_out_4_bits_fpWen),
    .io_out_4_bits_vecWen(io_out_4_bits_vecWen),
    .io_out_4_bits_v0Wen(io_out_4_bits_v0Wen),
    .io_out_4_bits_vlWen(io_out_4_bits_vlWen),
    .io_out_4_bits_isXSTrap(io_out_4_bits_isXSTrap),
    .io_out_4_bits_waitForward(io_out_4_bits_waitForward),
    .io_out_4_bits_blockBackward(io_out_4_bits_blockBackward),
    .io_out_4_bits_flushPipe(io_out_4_bits_flushPipe),
    .io_out_4_bits_canRobCompress(io_out_4_bits_canRobCompress),
    .io_out_4_bits_selImm(io_out_4_bits_selImm),
    .io_out_4_bits_imm(io_out_4_bits_imm),
    .io_out_4_bits_fpu_typeTagOut(io_out_4_bits_fpu_typeTagOut),
    .io_out_4_bits_fpu_wflags(io_out_4_bits_fpu_wflags),
    .io_out_4_bits_fpu_typ(io_out_4_bits_fpu_typ),
    .io_out_4_bits_fpu_fmt(io_out_4_bits_fpu_fmt),
    .io_out_4_bits_fpu_rm(io_out_4_bits_fpu_rm),
    .io_out_4_bits_vpu_vill(io_out_4_bits_vpu_vill),
    .io_out_4_bits_vpu_vma(io_out_4_bits_vpu_vma),
    .io_out_4_bits_vpu_vta(io_out_4_bits_vpu_vta),
    .io_out_4_bits_vpu_vsew(io_out_4_bits_vpu_vsew),
    .io_out_4_bits_vpu_vlmul(io_out_4_bits_vpu_vlmul),
    .io_out_4_bits_vpu_specVill(io_out_4_bits_vpu_specVill),
    .io_out_4_bits_vpu_specVma(io_out_4_bits_vpu_specVma),
    .io_out_4_bits_vpu_specVta(io_out_4_bits_vpu_specVta),
    .io_out_4_bits_vpu_specVsew(io_out_4_bits_vpu_specVsew),
    .io_out_4_bits_vpu_specVlmul(io_out_4_bits_vpu_specVlmul),
    .io_out_4_bits_vpu_vm(io_out_4_bits_vpu_vm),
    .io_out_4_bits_vpu_vstart(io_out_4_bits_vpu_vstart),
    .io_out_4_bits_vpu_fpu_isFoldTo1_2(io_out_4_bits_vpu_fpu_isFoldTo1_2),
    .io_out_4_bits_vpu_fpu_isFoldTo1_4(io_out_4_bits_vpu_fpu_isFoldTo1_4),
    .io_out_4_bits_vpu_fpu_isFoldTo1_8(io_out_4_bits_vpu_fpu_isFoldTo1_8),
    .io_out_4_bits_vpu_nf(io_out_4_bits_vpu_nf),
    .io_out_4_bits_vpu_veew(io_out_4_bits_vpu_veew),
    .io_out_4_bits_vpu_isExt(io_out_4_bits_vpu_isExt),
    .io_out_4_bits_vpu_isNarrow(io_out_4_bits_vpu_isNarrow),
    .io_out_4_bits_vpu_isDstMask(io_out_4_bits_vpu_isDstMask),
    .io_out_4_bits_vpu_isOpMask(io_out_4_bits_vpu_isOpMask),
    .io_out_4_bits_vpu_isDependOldVd(io_out_4_bits_vpu_isDependOldVd),
    .io_out_4_bits_vpu_isWritePartVd(io_out_4_bits_vpu_isWritePartVd),
    .io_out_4_bits_vpu_isVleff(io_out_4_bits_vpu_isVleff),
    .io_out_4_bits_vlsInstr(io_out_4_bits_vlsInstr),
    .io_out_4_bits_wfflags(io_out_4_bits_wfflags),
    .io_out_4_bits_isMove(io_out_4_bits_isMove),
    .io_out_4_bits_uopIdx(io_out_4_bits_uopIdx),
    .io_out_4_bits_uopSplitType(io_out_4_bits_uopSplitType),
    .io_out_4_bits_isVset(io_out_4_bits_isVset),
    .io_out_4_bits_firstUop(io_out_4_bits_firstUop),
    .io_out_4_bits_lastUop(io_out_4_bits_lastUop),
    .io_out_4_bits_numWB(io_out_4_bits_numWB),
    .io_out_4_bits_commitType(io_out_4_bits_commitType),
    .io_out_5_ready(io_out_5_ready),
    .io_out_5_valid(io_out_5_valid),
    .io_out_5_bits_instr(io_out_5_bits_instr),
    .io_out_5_bits_exceptionVec_0(io_out_5_bits_exceptionVec_0),
    .io_out_5_bits_exceptionVec_1(io_out_5_bits_exceptionVec_1),
    .io_out_5_bits_exceptionVec_2(io_out_5_bits_exceptionVec_2),
    .io_out_5_bits_exceptionVec_3(io_out_5_bits_exceptionVec_3),
    .io_out_5_bits_exceptionVec_4(io_out_5_bits_exceptionVec_4),
    .io_out_5_bits_exceptionVec_5(io_out_5_bits_exceptionVec_5),
    .io_out_5_bits_exceptionVec_6(io_out_5_bits_exceptionVec_6),
    .io_out_5_bits_exceptionVec_7(io_out_5_bits_exceptionVec_7),
    .io_out_5_bits_exceptionVec_8(io_out_5_bits_exceptionVec_8),
    .io_out_5_bits_exceptionVec_9(io_out_5_bits_exceptionVec_9),
    .io_out_5_bits_exceptionVec_10(io_out_5_bits_exceptionVec_10),
    .io_out_5_bits_exceptionVec_11(io_out_5_bits_exceptionVec_11),
    .io_out_5_bits_exceptionVec_12(io_out_5_bits_exceptionVec_12),
    .io_out_5_bits_exceptionVec_13(io_out_5_bits_exceptionVec_13),
    .io_out_5_bits_exceptionVec_14(io_out_5_bits_exceptionVec_14),
    .io_out_5_bits_exceptionVec_15(io_out_5_bits_exceptionVec_15),
    .io_out_5_bits_exceptionVec_16(io_out_5_bits_exceptionVec_16),
    .io_out_5_bits_exceptionVec_17(io_out_5_bits_exceptionVec_17),
    .io_out_5_bits_exceptionVec_18(io_out_5_bits_exceptionVec_18),
    .io_out_5_bits_exceptionVec_19(io_out_5_bits_exceptionVec_19),
    .io_out_5_bits_exceptionVec_20(io_out_5_bits_exceptionVec_20),
    .io_out_5_bits_exceptionVec_21(io_out_5_bits_exceptionVec_21),
    .io_out_5_bits_exceptionVec_22(io_out_5_bits_exceptionVec_22),
    .io_out_5_bits_exceptionVec_23(io_out_5_bits_exceptionVec_23),
    .io_out_5_bits_isFetchMalAddr(io_out_5_bits_isFetchMalAddr),
    .io_out_5_bits_trigger(io_out_5_bits_trigger),
    .io_out_5_bits_preDecodeInfo_isRVC(io_out_5_bits_preDecodeInfo_isRVC),
    .io_out_5_bits_preDecodeInfo_brType(io_out_5_bits_preDecodeInfo_brType),
    .io_out_5_bits_pred_taken(io_out_5_bits_pred_taken),
    .io_out_5_bits_crossPageIPFFix(io_out_5_bits_crossPageIPFFix),
    .io_out_5_bits_ftqPtr_flag(io_out_5_bits_ftqPtr_flag),
    .io_out_5_bits_ftqPtr_value(io_out_5_bits_ftqPtr_value),
    .io_out_5_bits_ftqOffset(io_out_5_bits_ftqOffset),
    .io_out_5_bits_srcType_0(io_out_5_bits_srcType_0),
    .io_out_5_bits_srcType_1(io_out_5_bits_srcType_1),
    .io_out_5_bits_srcType_2(io_out_5_bits_srcType_2),
    .io_out_5_bits_srcType_3(io_out_5_bits_srcType_3),
    .io_out_5_bits_srcType_4(io_out_5_bits_srcType_4),
    .io_out_5_bits_lsrc_0(io_out_5_bits_lsrc_0),
    .io_out_5_bits_lsrc_1(io_out_5_bits_lsrc_1),
    .io_out_5_bits_lsrc_2(io_out_5_bits_lsrc_2),
    .io_out_5_bits_ldest(io_out_5_bits_ldest),
    .io_out_5_bits_fuType(io_out_5_bits_fuType),
    .io_out_5_bits_fuOpType(io_out_5_bits_fuOpType),
    .io_out_5_bits_rfWen(io_out_5_bits_rfWen),
    .io_out_5_bits_fpWen(io_out_5_bits_fpWen),
    .io_out_5_bits_vecWen(io_out_5_bits_vecWen),
    .io_out_5_bits_v0Wen(io_out_5_bits_v0Wen),
    .io_out_5_bits_vlWen(io_out_5_bits_vlWen),
    .io_out_5_bits_isXSTrap(io_out_5_bits_isXSTrap),
    .io_out_5_bits_waitForward(io_out_5_bits_waitForward),
    .io_out_5_bits_blockBackward(io_out_5_bits_blockBackward),
    .io_out_5_bits_flushPipe(io_out_5_bits_flushPipe),
    .io_out_5_bits_canRobCompress(io_out_5_bits_canRobCompress),
    .io_out_5_bits_selImm(io_out_5_bits_selImm),
    .io_out_5_bits_imm(io_out_5_bits_imm),
    .io_out_5_bits_fpu_typeTagOut(io_out_5_bits_fpu_typeTagOut),
    .io_out_5_bits_fpu_wflags(io_out_5_bits_fpu_wflags),
    .io_out_5_bits_fpu_typ(io_out_5_bits_fpu_typ),
    .io_out_5_bits_fpu_fmt(io_out_5_bits_fpu_fmt),
    .io_out_5_bits_fpu_rm(io_out_5_bits_fpu_rm),
    .io_out_5_bits_vpu_vill(io_out_5_bits_vpu_vill),
    .io_out_5_bits_vpu_vma(io_out_5_bits_vpu_vma),
    .io_out_5_bits_vpu_vta(io_out_5_bits_vpu_vta),
    .io_out_5_bits_vpu_vsew(io_out_5_bits_vpu_vsew),
    .io_out_5_bits_vpu_vlmul(io_out_5_bits_vpu_vlmul),
    .io_out_5_bits_vpu_specVill(io_out_5_bits_vpu_specVill),
    .io_out_5_bits_vpu_specVma(io_out_5_bits_vpu_specVma),
    .io_out_5_bits_vpu_specVta(io_out_5_bits_vpu_specVta),
    .io_out_5_bits_vpu_specVsew(io_out_5_bits_vpu_specVsew),
    .io_out_5_bits_vpu_specVlmul(io_out_5_bits_vpu_specVlmul),
    .io_out_5_bits_vpu_vm(io_out_5_bits_vpu_vm),
    .io_out_5_bits_vpu_vstart(io_out_5_bits_vpu_vstart),
    .io_out_5_bits_vpu_fpu_isFoldTo1_2(io_out_5_bits_vpu_fpu_isFoldTo1_2),
    .io_out_5_bits_vpu_fpu_isFoldTo1_4(io_out_5_bits_vpu_fpu_isFoldTo1_4),
    .io_out_5_bits_vpu_fpu_isFoldTo1_8(io_out_5_bits_vpu_fpu_isFoldTo1_8),
    .io_out_5_bits_vpu_nf(io_out_5_bits_vpu_nf),
    .io_out_5_bits_vpu_veew(io_out_5_bits_vpu_veew),
    .io_out_5_bits_vpu_isExt(io_out_5_bits_vpu_isExt),
    .io_out_5_bits_vpu_isNarrow(io_out_5_bits_vpu_isNarrow),
    .io_out_5_bits_vpu_isDstMask(io_out_5_bits_vpu_isDstMask),
    .io_out_5_bits_vpu_isOpMask(io_out_5_bits_vpu_isOpMask),
    .io_out_5_bits_vpu_isDependOldVd(io_out_5_bits_vpu_isDependOldVd),
    .io_out_5_bits_vpu_isWritePartVd(io_out_5_bits_vpu_isWritePartVd),
    .io_out_5_bits_vpu_isVleff(io_out_5_bits_vpu_isVleff),
    .io_out_5_bits_vlsInstr(io_out_5_bits_vlsInstr),
    .io_out_5_bits_wfflags(io_out_5_bits_wfflags),
    .io_out_5_bits_isMove(io_out_5_bits_isMove),
    .io_out_5_bits_uopIdx(io_out_5_bits_uopIdx),
    .io_out_5_bits_uopSplitType(io_out_5_bits_uopSplitType),
    .io_out_5_bits_isVset(io_out_5_bits_isVset),
    .io_out_5_bits_firstUop(io_out_5_bits_firstUop),
    .io_out_5_bits_lastUop(io_out_5_bits_lastUop),
    .io_out_5_bits_numWB(io_out_5_bits_numWB),
    .io_out_5_bits_commitType(io_out_5_bits_commitType),
    .io_intRat_0_0_hold(io_intRat_0_0_hold),
    .io_intRat_0_0_addr(io_intRat_0_0_addr),
    .io_intRat_0_1_hold(io_intRat_0_1_hold),
    .io_intRat_0_1_addr(io_intRat_0_1_addr),
    .io_intRat_1_0_hold(io_intRat_1_0_hold),
    .io_intRat_1_0_addr(io_intRat_1_0_addr),
    .io_intRat_1_1_hold(io_intRat_1_1_hold),
    .io_intRat_1_1_addr(io_intRat_1_1_addr),
    .io_intRat_2_0_hold(io_intRat_2_0_hold),
    .io_intRat_2_0_addr(io_intRat_2_0_addr),
    .io_intRat_2_1_hold(io_intRat_2_1_hold),
    .io_intRat_2_1_addr(io_intRat_2_1_addr),
    .io_intRat_3_0_hold(io_intRat_3_0_hold),
    .io_intRat_3_0_addr(io_intRat_3_0_addr),
    .io_intRat_3_1_hold(io_intRat_3_1_hold),
    .io_intRat_3_1_addr(io_intRat_3_1_addr),
    .io_intRat_4_0_hold(io_intRat_4_0_hold),
    .io_intRat_4_0_addr(io_intRat_4_0_addr),
    .io_intRat_4_1_hold(io_intRat_4_1_hold),
    .io_intRat_4_1_addr(io_intRat_4_1_addr),
    .io_intRat_5_0_hold(io_intRat_5_0_hold),
    .io_intRat_5_0_addr(io_intRat_5_0_addr),
    .io_intRat_5_1_hold(io_intRat_5_1_hold),
    .io_intRat_5_1_addr(io_intRat_5_1_addr),
    .io_fpRat_0_0_hold(io_fpRat_0_0_hold),
    .io_fpRat_0_0_addr(io_fpRat_0_0_addr),
    .io_fpRat_0_1_hold(io_fpRat_0_1_hold),
    .io_fpRat_0_1_addr(io_fpRat_0_1_addr),
    .io_fpRat_0_2_hold(io_fpRat_0_2_hold),
    .io_fpRat_0_2_addr(io_fpRat_0_2_addr),
    .io_fpRat_1_0_hold(io_fpRat_1_0_hold),
    .io_fpRat_1_0_addr(io_fpRat_1_0_addr),
    .io_fpRat_1_1_hold(io_fpRat_1_1_hold),
    .io_fpRat_1_1_addr(io_fpRat_1_1_addr),
    .io_fpRat_1_2_hold(io_fpRat_1_2_hold),
    .io_fpRat_1_2_addr(io_fpRat_1_2_addr),
    .io_fpRat_2_0_hold(io_fpRat_2_0_hold),
    .io_fpRat_2_0_addr(io_fpRat_2_0_addr),
    .io_fpRat_2_1_hold(io_fpRat_2_1_hold),
    .io_fpRat_2_1_addr(io_fpRat_2_1_addr),
    .io_fpRat_2_2_hold(io_fpRat_2_2_hold),
    .io_fpRat_2_2_addr(io_fpRat_2_2_addr),
    .io_fpRat_3_0_hold(io_fpRat_3_0_hold),
    .io_fpRat_3_0_addr(io_fpRat_3_0_addr),
    .io_fpRat_3_1_hold(io_fpRat_3_1_hold),
    .io_fpRat_3_1_addr(io_fpRat_3_1_addr),
    .io_fpRat_3_2_hold(io_fpRat_3_2_hold),
    .io_fpRat_3_2_addr(io_fpRat_3_2_addr),
    .io_fpRat_4_0_hold(io_fpRat_4_0_hold),
    .io_fpRat_4_0_addr(io_fpRat_4_0_addr),
    .io_fpRat_4_1_hold(io_fpRat_4_1_hold),
    .io_fpRat_4_1_addr(io_fpRat_4_1_addr),
    .io_fpRat_4_2_hold(io_fpRat_4_2_hold),
    .io_fpRat_4_2_addr(io_fpRat_4_2_addr),
    .io_fpRat_5_0_hold(io_fpRat_5_0_hold),
    .io_fpRat_5_0_addr(io_fpRat_5_0_addr),
    .io_fpRat_5_1_hold(io_fpRat_5_1_hold),
    .io_fpRat_5_1_addr(io_fpRat_5_1_addr),
    .io_fpRat_5_2_hold(io_fpRat_5_2_hold),
    .io_fpRat_5_2_addr(io_fpRat_5_2_addr),
    .io_vecRat_0_0_hold(io_vecRat_0_0_hold),
    .io_vecRat_0_0_addr(io_vecRat_0_0_addr),
    .io_vecRat_0_1_hold(io_vecRat_0_1_hold),
    .io_vecRat_0_1_addr(io_vecRat_0_1_addr),
    .io_vecRat_0_2_hold(io_vecRat_0_2_hold),
    .io_vecRat_0_2_addr(io_vecRat_0_2_addr),
    .io_vecRat_1_0_hold(io_vecRat_1_0_hold),
    .io_vecRat_1_0_addr(io_vecRat_1_0_addr),
    .io_vecRat_1_1_hold(io_vecRat_1_1_hold),
    .io_vecRat_1_1_addr(io_vecRat_1_1_addr),
    .io_vecRat_1_2_hold(io_vecRat_1_2_hold),
    .io_vecRat_1_2_addr(io_vecRat_1_2_addr),
    .io_vecRat_2_0_hold(io_vecRat_2_0_hold),
    .io_vecRat_2_0_addr(io_vecRat_2_0_addr),
    .io_vecRat_2_1_hold(io_vecRat_2_1_hold),
    .io_vecRat_2_1_addr(io_vecRat_2_1_addr),
    .io_vecRat_2_2_hold(io_vecRat_2_2_hold),
    .io_vecRat_2_2_addr(io_vecRat_2_2_addr),
    .io_vecRat_3_0_hold(io_vecRat_3_0_hold),
    .io_vecRat_3_0_addr(io_vecRat_3_0_addr),
    .io_vecRat_3_1_hold(io_vecRat_3_1_hold),
    .io_vecRat_3_1_addr(io_vecRat_3_1_addr),
    .io_vecRat_3_2_hold(io_vecRat_3_2_hold),
    .io_vecRat_3_2_addr(io_vecRat_3_2_addr),
    .io_vecRat_4_0_hold(io_vecRat_4_0_hold),
    .io_vecRat_4_0_addr(io_vecRat_4_0_addr),
    .io_vecRat_4_1_hold(io_vecRat_4_1_hold),
    .io_vecRat_4_1_addr(io_vecRat_4_1_addr),
    .io_vecRat_4_2_hold(io_vecRat_4_2_hold),
    .io_vecRat_4_2_addr(io_vecRat_4_2_addr),
    .io_vecRat_5_0_hold(io_vecRat_5_0_hold),
    .io_vecRat_5_0_addr(io_vecRat_5_0_addr),
    .io_vecRat_5_1_hold(io_vecRat_5_1_hold),
    .io_vecRat_5_1_addr(io_vecRat_5_1_addr),
    .io_vecRat_5_2_hold(io_vecRat_5_2_hold),
    .io_vecRat_5_2_addr(io_vecRat_5_2_addr),
    .io_csrCtrl_singlestep(io_csrCtrl_singlestep),
    .io_fromCSR_illegalInst_sfenceVMA(io_fromCSR_illegalInst_sfenceVMA),
    .io_fromCSR_illegalInst_sfencePart(io_fromCSR_illegalInst_sfencePart),
    .io_fromCSR_illegalInst_hfenceGVMA(io_fromCSR_illegalInst_hfenceGVMA),
    .io_fromCSR_illegalInst_hfenceVVMA(io_fromCSR_illegalInst_hfenceVVMA),
    .io_fromCSR_illegalInst_hlsv(io_fromCSR_illegalInst_hlsv),
    .io_fromCSR_illegalInst_fsIsOff(io_fromCSR_illegalInst_fsIsOff),
    .io_fromCSR_illegalInst_vsIsOff(io_fromCSR_illegalInst_vsIsOff),
    .io_fromCSR_illegalInst_wfi(io_fromCSR_illegalInst_wfi),
    .io_fromCSR_illegalInst_frm(io_fromCSR_illegalInst_frm),
    .io_fromCSR_illegalInst_cboZ(io_fromCSR_illegalInst_cboZ),
    .io_fromCSR_illegalInst_cboCF(io_fromCSR_illegalInst_cboCF),
    .io_fromCSR_illegalInst_cboI(io_fromCSR_illegalInst_cboI),
    .io_fromCSR_virtualInst_sfenceVMA(io_fromCSR_virtualInst_sfenceVMA),
    .io_fromCSR_virtualInst_sfencePart(io_fromCSR_virtualInst_sfencePart),
    .io_fromCSR_virtualInst_hfence(io_fromCSR_virtualInst_hfence),
    .io_fromCSR_virtualInst_hlsv(io_fromCSR_virtualInst_hlsv),
    .io_fromCSR_virtualInst_wfi(io_fromCSR_virtualInst_wfi),
    .io_fromCSR_virtualInst_cboZ(io_fromCSR_virtualInst_cboZ),
    .io_fromCSR_virtualInst_cboCF(io_fromCSR_virtualInst_cboCF),
    .io_fromCSR_virtualInst_cboI(io_fromCSR_virtualInst_cboI),
    .io_fromCSR_special_cboI2F(io_fromCSR_special_cboI2F),
    .io_fusion_0(io_fusion_0),
    .io_fusion_1(io_fusion_1),
    .io_fusion_2(io_fusion_2),
    .io_fusion_3(io_fusion_3),
    .io_fusion_4(io_fusion_4),
    .io_fromRob_isResumeVType(io_fromRob_isResumeVType),
    .io_fromRob_walkToArchVType(io_fromRob_walkToArchVType),
    .io_fromRob_commitVType_vtype_valid(io_fromRob_commitVType_vtype_valid),
    .io_fromRob_commitVType_vtype_bits_illegal(io_fromRob_commitVType_vtype_bits_illegal),
    .io_fromRob_commitVType_vtype_bits_vma(io_fromRob_commitVType_vtype_bits_vma),
    .io_fromRob_commitVType_vtype_bits_vta(io_fromRob_commitVType_vtype_bits_vta),
    .io_fromRob_commitVType_vtype_bits_vsew(io_fromRob_commitVType_vtype_bits_vsew),
    .io_fromRob_commitVType_vtype_bits_vlmul(io_fromRob_commitVType_vtype_bits_vlmul),
    .io_fromRob_commitVType_hasVsetvl(io_fromRob_commitVType_hasVsetvl),
    .io_fromRob_walkVType_valid(io_fromRob_walkVType_valid),
    .io_fromRob_walkVType_bits_illegal(io_fromRob_walkVType_bits_illegal),
    .io_fromRob_walkVType_bits_vma(io_fromRob_walkVType_bits_vma),
    .io_fromRob_walkVType_bits_vta(io_fromRob_walkVType_bits_vta),
    .io_fromRob_walkVType_bits_vsew(io_fromRob_walkVType_bits_vsew),
    .io_fromRob_walkVType_bits_vlmul(io_fromRob_walkVType_bits_vlmul),
    .io_vsetvlVType_illegal(io_vsetvlVType_illegal),
    .io_vsetvlVType_vma(io_vsetvlVType_vma),
    .io_vsetvlVType_vta(io_vsetvlVType_vta),
    .io_vsetvlVType_vsew(io_vsetvlVType_vsew),
    .io_vsetvlVType_vlmul(io_vsetvlVType_vlmul),
    .io_vstart(io_vstart),
    .io_toCSR_trapInstInfo_valid(io_toCSR_trapInstInfo_valid),
    .io_toCSR_trapInstInfo_bits_instr(io_toCSR_trapInstInfo_bits_instr),
    .io_toCSR_trapInstInfo_bits_ftqPtr_flag(io_toCSR_trapInstInfo_bits_ftqPtr_flag),
    .io_toCSR_trapInstInfo_bits_ftqPtr_value(io_toCSR_trapInstInfo_bits_ftqPtr_value),
    .io_toCSR_trapInstInfo_bits_ftqOffset(io_toCSR_trapInstInfo_bits_ftqOffset),
    .io_perf_0_value(io_perf_0_value),
    .io_perf_1_value(io_perf_1_value),
    .io_perf_2_value(io_perf_2_value),
    .io_perf_3_value(io_perf_3_value)
 );


endmodule
